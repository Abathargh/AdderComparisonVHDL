library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TB_RCA is
    generic(width: integer := 16);
end TB_RCA;

architecture Behavioral of TB_RCA is

component RCA_3IN
    Port(
        A, B, C: in std_logic_vector(width - 1 downto 0);
        clk: in std_logic;
        Sum: out std_logic_vector(width + 1 downto 0)
    );
end component;

signal A, B, C: std_logic_vector(width - 1 downto 0);
signal clk: std_logic;
signal Sum: std_logic_vector(width + 1 downto 0);

constant clk_period : time := 3 ns;

begin
    uut: RCA_3IN port map(A => A, B => B, C => C, clk => clk, Sum => Sum);
    
    process begin
        clk <= '0';
        wait for clk_period / 2;
        clk <= '1';
        wait for clk_period / 2;
    end process;
    
    process begin
        wait for 100 ns;
        A <= "1110111010100100";
        B <= "0111000011101101";
        C <= "1111011111101010";
        wait for clk_period;
        A <= "1011100000110001";
        B <= "1111100110011000";
        C <= "1100010000101000";
        wait for clk_period;
        A <= "1101010011100010";
        B <= "1000011011110111";
        C <= "0111111010010000";
        wait for clk_period;
        A <= "1100011110110101";
        B <= "1000110000100001";
        C <= "0000010111111011";
        wait for clk_period;
        A <= "1111011001101011";
        B <= "0011110000100100";
        C <= "0111000111101001";
        wait for clk_period;
        A <= "0001001001110000";
        B <= "0110101010011110";
        C <= "0111011000100111";
        wait for clk_period;
        A <= "0101011011110101";
        B <= "1011010101110001";
        C <= "0110000111010010";
        wait for clk_period;
        A <= "1011011010111011";
        B <= "0000001010100100";
        C <= "0111011010111101";
        wait for clk_period;
        A <= "1110000100101100";
        B <= "0101111001010010";
        C <= "0100100010100000";
        wait for clk_period;
        A <= "0111110011001010";
        B <= "1000010100100001";
        C <= "0000001111101011";
        wait for clk_period;
        A <= "0001000111011110";
        B <= "0010100100010100";
        C <= "1101011101110100";
        wait for clk_period;
        A <= "1011111011001101";
        B <= "0111011100100001";
        C <= "1001001011010101";
        wait for clk_period;
        A <= "1010010011110011";
        B <= "1111011011110000";
        C <= "1110101001101011";
        wait for clk_period;
        A <= "1110100111001111";
        B <= "1101000000110011";
        C <= "1001001000000110";
        wait for clk_period;
        A <= "1100110101101011";
        B <= "1101010000100110";
        C <= "0000101111110011";
        wait for clk_period;
        A <= "0011010110111101";
        B <= "0000010110110100";
        C <= "1111100100001101";
        wait for clk_period;
        A <= "1000010101101111";
        B <= "0011110110111100";
        C <= "1101110110000111";
        wait for clk_period;
        A <= "1111010110010001";
        B <= "1000011101001111";
        C <= "1100111011001000";
        wait for clk_period;
        A <= "0001011000011111";
        B <= "0011100100100111";
        C <= "0111101000111101";
        wait for clk_period;
        A <= "1010101110010111";
        B <= "0111111111011010";
        C <= "1110110110000000";
        wait for clk_period;
        A <= "0000010111010100";
        B <= "0001101100101100";
        C <= "0010010001101010";
        wait for clk_period;
        A <= "1001101111111001";
        B <= "1100101011110111";
        C <= "0010101010000010";
        wait for clk_period;
        A <= "1111110011011101";
        B <= "1111000111111000";
        C <= "0110010011000111";
        wait for clk_period;
        A <= "1111000001101010";
        B <= "1110100000010010";
        C <= "0010010110110010";
        wait for clk_period;
        A <= "0000001100011110";
        B <= "0101100101001000";
        C <= "1111100111011100";
        wait for clk_period;
        A <= "0111101111110110";
        B <= "0110101010101110";
        C <= "0101000011010100";
        wait for clk_period;
        A <= "1100010001111101";
        B <= "1111101101011010";
        C <= "0010100110101010";
        wait for clk_period;
        A <= "1111111001000010";
        B <= "1110011000100010";
        C <= "0000011101111000";
        wait for clk_period;
        A <= "0110001011100000";
        B <= "1000001001100010";
        C <= "1011101011011010";
        wait for clk_period;
        A <= "1100010010110000";
        B <= "1111111001110101";
        C <= "1111000011110110";
        wait for clk_period;
        A <= "0110110001001110";
        B <= "1101000001101010";
        C <= "1110010101010100";
        wait for clk_period;
        A <= "1010010101000000";
        B <= "0011111101101011";
        C <= "0110100011111011";
        wait for clk_period;
        A <= "1110100111111000";
        B <= "1110010011011110";
        C <= "1010001101010010";
        wait for clk_period;
        A <= "1010110010011110";
        B <= "0001101011000111";
        C <= "1011100100111101";
        wait for clk_period;
        A <= "1011001101101011";
        B <= "1011110111101001";
        C <= "0000111100010100";
        wait for clk_period;
        A <= "1010010011001101";
        B <= "1111110101010001";
        C <= "0110001000101010";
        wait for clk_period;
        A <= "1000100000111110";
        B <= "0000010100101100";
        C <= "0111010010111001";
        wait for clk_period;
        A <= "1001100010101110";
        B <= "0110101111000010";
        C <= "1111100000011111";
        wait for clk_period;
        A <= "1010011100110100";
        B <= "0011011011111110";
        C <= "0000110111101100";
        wait for clk_period;
        A <= "1010011101010000";
        B <= "0011001100011110";
        C <= "0101100010001100";
        wait for clk_period;
        A <= "1101111111101111";
        B <= "0100001100000000";
        C <= "0000110011100011";
        wait for clk_period;
        A <= "1110101101100101";
        B <= "0110010100111001";
        C <= "1111111100011100";
        wait for clk_period;
        A <= "1110001010111111";
        B <= "1110100011001111";
        C <= "1110100001111111";
        wait for clk_period;
        A <= "1010000011011101";
        B <= "0111110000100111";
        C <= "1110100101011001";
        wait for clk_period;
        A <= "1010100111001001";
        B <= "1000111000000110";
        C <= "1011111101010110";
        wait for clk_period;
        A <= "0010100101011110";
        B <= "1000011101111101";
        C <= "0111100010111111";
        wait for clk_period;
        A <= "0101111110110011";
        B <= "0101101110110111";
        C <= "1100011011101001";
        wait for clk_period;
        A <= "0110111110010111";
        B <= "0010100110111101";
        C <= "0010001000100000";
        wait for clk_period;
        A <= "1101110100000011";
        B <= "1100000000001111";
        C <= "1101110101100001";
        wait for clk_period;
        A <= "1111010001101000";
        B <= "1011010110111110";
        C <= "1010001000101110";
        wait for clk_period;
        A <= "0101010110100101";
        B <= "1000011100011100";
        C <= "1110011110100010";
        wait for clk_period;
        A <= "0000101101110011";
        B <= "1011011001110101";
        C <= "0001111000011000";
        wait for clk_period;
        A <= "0101111100000111";
        B <= "0011111110000110";
        C <= "0011010100001111";
        wait for clk_period;
        A <= "0011011011011101";
        B <= "0001101001000001";
        C <= "1100110010101111";
        wait for clk_period;
        A <= "0010101101110001";
        B <= "0010101010101011";
        C <= "1000011110111110";
        wait for clk_period;
        A <= "1001011100110111";
        B <= "0011100111010010";
        C <= "0100001001111000";
        wait for clk_period;
        A <= "1111011100110111";
        B <= "1100100010111100";
        C <= "0100001110001011";
        wait for clk_period;
        A <= "1111101001100111";
        B <= "0100111001001100";
        C <= "0110001110111110";
        wait for clk_period;
        A <= "0000110101000011";
        B <= "0011010001001110";
        C <= "1100101010010010";
        wait for clk_period;
        A <= "1011111001010111";
        B <= "1010001100000010";
        C <= "1000110101110011";
        wait for clk_period;
        A <= "1111110011011110";
        B <= "1010001100101010";
        C <= "1001011000011001";
        wait for clk_period;
        A <= "1001110010100101";
        B <= "1101100000100010";
        C <= "0000010101111110";
        wait for clk_period;
        A <= "0101010110100010";
        B <= "1110100111101010";
        C <= "0001100100000111";
        wait for clk_period;
        A <= "1110000010001001";
        B <= "0100111011011010";
        C <= "1100101010000001";
        wait for clk_period;
        A <= "0011011000010010";
        B <= "0101011000111010";
        C <= "1100100111011101";
        wait for clk_period;
        A <= "1001110001000001";
        B <= "1101001001010000";
        C <= "0001010011010110";
        wait for clk_period;
        A <= "1100010111110101";
        B <= "1100011010010011";
        C <= "0101101010111101";
        wait for clk_period;
        A <= "1111000001111011";
        B <= "1000001110000111";
        C <= "0101001110000111";
        wait for clk_period;
        A <= "1110100011010010";
        B <= "0110001111000100";
        C <= "0110110110001000";
        wait for clk_period;
        A <= "1010000110010110";
        B <= "0000100011110000";
        C <= "0011000011111010";
        wait for clk_period;
        A <= "0111111111111100";
        B <= "1101110010000011";
        C <= "1100110000010101";
        wait for clk_period;
        A <= "0110101001000110";
        B <= "1101011001001110";
        C <= "0011101100010011";
        wait for clk_period;
        A <= "1001011110101001";
        B <= "0111110111000100";
        C <= "1110100000011010";
        wait for clk_period;
        A <= "0111011001111100";
        B <= "0001100001111110";
        C <= "1000010000010010";
        wait for clk_period;
        A <= "1101011010001111";
        B <= "1011110000100100";
        C <= "0111010111001111";
        wait for clk_period;
        A <= "0101010011111110";
        B <= "0001111000101010";
        C <= "0111101001011110";
        wait for clk_period;
        A <= "0100001011111000";
        B <= "1001010010011101";
        C <= "0110010100101011";
        wait for clk_period;
        A <= "1111001000100111";
        B <= "0111011011101101";
        C <= "1100101100000001";
        wait for clk_period;
        A <= "0111011101110001";
        B <= "1000010111101001";
        C <= "1011110011000010";
        wait for clk_period;
        A <= "1110100101111101";
        B <= "0101011101100110";
        C <= "0011100111010110";
        wait for clk_period;
        A <= "0000011111011110";
        B <= "0000011010000000";
        C <= "0111111000101101";
        wait for clk_period;
        A <= "1101111110110110";
        B <= "0000101001000101";
        C <= "1011100111111111";
        wait for clk_period;
        A <= "0011000110111111";
        B <= "1110101101010100";
        C <= "1111101101011100";
        wait for clk_period;
        A <= "1000111001011011";
        B <= "1110011111010011";
        C <= "0111001001101111";
        wait for clk_period;
        A <= "1001101000110000";
        B <= "1001010100100101";
        C <= "0011100011010110";
        wait for clk_period;
        A <= "0101111011011000";
        B <= "0101011100010101";
        C <= "1000011001110100";
        wait for clk_period;
        A <= "1001011000001110";
        B <= "1011101011110001";
        C <= "0100100111011001";
        wait for clk_period;
        A <= "1100110011100001";
        B <= "0101000011000010";
        C <= "0010100011010111";
        wait for clk_period;
        A <= "0011011100001000";
        B <= "1101010011000010";
        C <= "0011111000100101";
        wait for clk_period;
        A <= "0111110000011010";
        B <= "1001000011011000";
        C <= "1010000111010000";
        wait for clk_period;
        A <= "0111000001101010";
        B <= "0011101111011010";
        C <= "1000001111111110";
        wait for clk_period;
        A <= "0010000000110100";
        B <= "0011111000101111";
        C <= "0100110001101101";
        wait for clk_period;
        A <= "0111111101011111";
        B <= "1011111110000110";
        C <= "1000001100101000";
        wait for clk_period;
        A <= "1110110010111111";
        B <= "0011011101010111";
        C <= "1111110110110011";
        wait for clk_period;
        A <= "0011111011011111";
        B <= "1011100100000110";
        C <= "0100100110001100";
        wait for clk_period;
        A <= "0000000000101011";
        B <= "0000110010100111";
        C <= "1111100101110011";
        wait for clk_period;
        A <= "1100001110111010";
        B <= "1001111000000011";
        C <= "0100000101001111";
        wait for clk_period;
        A <= "0100101100111001";
        B <= "1011000100000111";
        C <= "0010011111101110";
        wait for clk_period;
        A <= "0011101001100010";
        B <= "1110011110110011";
        C <= "0111100001110100";
        wait for clk_period;
        A <= "0000101000100111";
        B <= "1100000001101001";
        C <= "1111101010101110";
        wait for clk_period;
        A <= "1011011101011001";
        B <= "1001111000001110";
        C <= "1011000101000011";
        wait for clk_period;
        A <= "1111101101011000";
        B <= "0110110110011010";
        C <= "0010111110111110";
        wait for clk_period;
        A <= "1001011001001100";
        B <= "1100001100010101";
        C <= "0001010101011000";
        wait for clk_period;
        A <= "1000001000100011";
        B <= "0011010011100000";
        C <= "0100000000010111";
        wait for clk_period;
        A <= "0001010010010111";
        B <= "0011011011000101";
        C <= "0110100100000011";
        wait for clk_period;
        A <= "1101010100111001";
        B <= "1110101111111010";
        C <= "1110101000110011";
        wait for clk_period;
        A <= "1010010100000111";
        B <= "0100001101110101";
        C <= "0010011110100111";
        wait for clk_period;
        A <= "0010001111100110";
        B <= "0000110000101011";
        C <= "0000001010100110";
        wait for clk_period;
        A <= "0101110000111001";
        B <= "1010100111110001";
        C <= "1000100100101100";
        wait for clk_period;
        A <= "0001000010100100";
        B <= "0001010100010000";
        C <= "0101010010110010";
        wait for clk_period;
        A <= "0101101111111010";
        B <= "1011010101000111";
        C <= "0010011011000010";
        wait for clk_period;
        A <= "0011010100011010";
        B <= "1110000010110110";
        C <= "0000000000111111";
        wait for clk_period;
        A <= "0101110110000111";
        B <= "1001011010111101";
        C <= "0011011101101101";
        wait for clk_period;
        A <= "0101010111001101";
        B <= "0110000110001011";
        C <= "0110111010011000";
        wait for clk_period;
        A <= "0110110011101111";
        B <= "1101111110100111";
        C <= "0110011111010001";
        wait for clk_period;
        A <= "1111110010100100";
        B <= "0001001100010100";
        C <= "0001011001111001";
        wait for clk_period;
        A <= "0100001100001011";
        B <= "0100111000100011";
        C <= "0100010110011011";
        wait for clk_period;
        A <= "1101001100000110";
        B <= "0010101001110011";
        C <= "1010000101101011";
        wait for clk_period;
        A <= "1010001010100000";
        B <= "0111000011110100";
        C <= "0010000100001011";
        wait for clk_period;
        A <= "1001111010001110";
        B <= "0010001011011100";
        C <= "1000101011101101";
        wait for clk_period;
        A <= "0110000010111001";
        B <= "1111001001010001";
        C <= "1100011010010101";
        wait for clk_period;
        A <= "1010110111111010";
        B <= "1111100011110100";
        C <= "0101110111001011";
        wait for clk_period;
        A <= "0010111010110000";
        B <= "0010000110001010";
        C <= "1110011000011111";
        wait for clk_period;
        A <= "0101100010011001";
        B <= "1011001010000101";
        C <= "1110110010110001";
        wait for clk_period;
        A <= "0111111110111100";
        B <= "1010100000111011";
        C <= "0110101111111100";
        wait for clk_period;
        A <= "0101100100111101";
        B <= "0100100101010000";
        C <= "0100010111011100";
        wait for clk_period;
        A <= "1100010011110010";
        B <= "1011101010110000";
        C <= "0001001000000011";
        wait for clk_period;
        A <= "0100100110100000";
        B <= "0010001101010011";
        C <= "1001111000111010";
        wait for clk_period;
        A <= "0000000010111110";
        B <= "1100001010000011";
        C <= "0100101011110010";
        wait for clk_period;
        A <= "0000000011100000";
        B <= "1000111010101111";
        C <= "0011000010011001";
        wait for clk_period;
        A <= "0001101000100101";
        B <= "0111110001101011";
        C <= "0010011100110000";
        wait for clk_period;
        A <= "1000001111011001";
        B <= "1101010010000001";
        C <= "1001010111001110";
        wait for clk_period;
        A <= "0010010010111000";
        B <= "0100001101001011";
        C <= "0010101011100110";
        wait for clk_period;
        A <= "1100010010110011";
        B <= "1111001011111110";
        C <= "0000100010100111";
        wait for clk_period;
        A <= "1001100101100110";
        B <= "1111110001100001";
        C <= "0011111001110010";
        wait for clk_period;
        A <= "1101111101100100";
        B <= "0101110001011010";
        C <= "1100110100100101";
        wait for clk_period;
        A <= "1010010010010000";
        B <= "0100000101100000";
        C <= "1101111110000110";
        wait for clk_period;
        A <= "0000101110000100";
        B <= "0010010001101000";
        C <= "1110110000011110";
        wait for clk_period;
        A <= "1101110101011101";
        B <= "0110010010011100";
        C <= "1110000100000010";
        wait for clk_period;
        A <= "0010010001101111";
        B <= "1110100011010111";
        C <= "0110110111000110";
        wait for clk_period;
        A <= "0100111010100000";
        B <= "0110010101110111";
        C <= "1111101100110101";
        wait for clk_period;
        A <= "0110100110010001";
        B <= "0110000110010011";
        C <= "0011010111110010";
        wait for clk_period;
        A <= "0010011100011010";
        B <= "0110101101111000";
        C <= "0101001101111101";
        wait for clk_period;
        A <= "1000101001111000";
        B <= "1100101000101011";
        C <= "1011110110111110";
        wait for clk_period;
        A <= "1100001011010101";
        B <= "1100100101111000";
        C <= "0110111101000111";
        wait for clk_period;
        A <= "1101010011100011";
        B <= "0001111011000011";
        C <= "0110110011110101";
        wait for clk_period;
        A <= "1111110001110010";
        B <= "1010001001110101";
        C <= "0111010101000101";
        wait for clk_period;
        A <= "0110100110001011";
        B <= "0111010000110000";
        C <= "0011010010111101";
        wait for clk_period;
        A <= "1010101010110110";
        B <= "0100011001001001";
        C <= "0010111110011111";
        wait for clk_period;
        A <= "1010001011010111";
        B <= "0110111101000010";
        C <= "0110000101000110";
        wait for clk_period;
        A <= "1000000000110110";
        B <= "0001100110010001";
        C <= "1101101011110100";
        wait for clk_period;
        A <= "0111000000001000";
        B <= "0001100011100001";
        C <= "0001110100100111";
        wait for clk_period;
        A <= "1111011010001001";
        B <= "0101100011111010";
        C <= "1101010100000011";
        wait for clk_period;
        A <= "0001100000100001";
        B <= "0111011001100000";
        C <= "1111000001010010";
        wait for clk_period;
        A <= "1000101000101110";
        B <= "0010100101101011";
        C <= "0011110000101101";
        wait for clk_period;
        A <= "1101100011000101";
        B <= "0010001001011110";
        C <= "0111110100100000";
        wait for clk_period;
        A <= "0011110101100000";
        B <= "1101010111111110";
        C <= "0100111110011010";
        wait for clk_period;
        A <= "1101111110010110";
        B <= "0110110100100011";
        C <= "0111111100010001";
        wait for clk_period;
        A <= "1101001100010100";
        B <= "1001011110110000";
        C <= "1100001001001100";
        wait for clk_period;
        A <= "0101000000100110";
        B <= "1100111101111000";
        C <= "0010100100010110";
        wait for clk_period;
        A <= "1001100010100100";
        B <= "1100011111111010";
        C <= "0010011101100011";
        wait for clk_period;
        A <= "1000100110101011";
        B <= "0001100100101101";
        C <= "1110000010111011";
        wait for clk_period;
        A <= "1100001000000000";
        B <= "0100110111001101";
        C <= "0011101011000100";
        wait for clk_period;
        A <= "1010010001011100";
        B <= "0001101100001011";
        C <= "1100000111101010";
        wait for clk_period;
        A <= "0110000011110100";
        B <= "1100011000001001";
        C <= "0010011000001101";
        wait for clk_period;
        A <= "0111110110101001";
        B <= "1100010001010010";
        C <= "1101001000110001";
        wait for clk_period;
        A <= "0010000011011001";
        B <= "0111000000001111";
        C <= "1000100101001001";
        wait for clk_period;
        A <= "0101110110001101";
        B <= "1100010010010000";
        C <= "0000000101001111";
        wait for clk_period;
        A <= "0010110010101101";
        B <= "0111100101110000";
        C <= "0010110011100010";
        wait for clk_period;
        A <= "1010111000100110";
        B <= "1010101010000000";
        C <= "0011101100111100";
        wait for clk_period;
        A <= "0110010010010110";
        B <= "0111111010111100";
        C <= "0100110100101000";
        wait for clk_period;
        A <= "0010010101010000";
        B <= "1000101010111001";
        C <= "0100001101110100";
        wait for clk_period;
        A <= "1100011101010111";
        B <= "0001000010010000";
        C <= "0010001100001110";
        wait for clk_period;
        A <= "1010001100000100";
        B <= "0000001000101011";
        C <= "1001110110101001";
        wait for clk_period;
        A <= "0001000000010000";
        B <= "0001000000000110";
        C <= "1000001101011001";
        wait for clk_period;
        A <= "0000110110101111";
        B <= "0110100001001001";
        C <= "0001110100011010";
        wait for clk_period;
        A <= "0101000010110111";
        B <= "1100000000101011";
        C <= "0110111110110111";
        wait for clk_period;
        A <= "0111000000001010";
        B <= "0000111111010101";
        C <= "0000011001001010";
        wait for clk_period;
        A <= "0110011010101011";
        B <= "1101000000001000";
        C <= "1001000000110011";
        wait for clk_period;
        A <= "0010100000010100";
        B <= "1100001110011110";
        C <= "0111010001001010";
        wait for clk_period;
        A <= "0000010101011101";
        B <= "1011011010100011";
        C <= "0001001011110100";
        wait for clk_period;
        A <= "0010011010010110";
        B <= "0111010000001010";
        C <= "0011001100010101";
        wait for clk_period;
        A <= "0011000101000010";
        B <= "0101010101111110";
        C <= "1110110100111001";
        wait for clk_period;
        A <= "1011011010111000";
        B <= "0101001100100010";
        C <= "1000000000011110";
        wait for clk_period;
        A <= "0100011101101101";
        B <= "0010110101100001";
        C <= "0101010000000010";
        wait for clk_period;
        A <= "1001111110001110";
        B <= "0011110000110010";
        C <= "0011011100110100";
        wait for clk_period;
        A <= "0101111001100010";
        B <= "1101010000110100";
        C <= "0011000011010100";
        wait for clk_period;
        A <= "1110010111011000";
        B <= "1011010010001000";
        C <= "0011011110000100";
        wait for clk_period;
        A <= "0011100000001011";
        B <= "0110100110110001";
        C <= "0101001100000001";
        wait for clk_period;
        A <= "1100111010111110";
        B <= "0010111011001101";
        C <= "1000000100111000";
        wait for clk_period;
        A <= "0010100000001110";
        B <= "1101111011111111";
        C <= "0110011010110010";
        wait for clk_period;
        A <= "1001111111100110";
        B <= "0010000100000000";
        C <= "0001000110011001";
        wait for clk_period;
        A <= "1111110100100101";
        B <= "1101101001101100";
        C <= "0100011111110001";
        wait for clk_period;
        A <= "0011110011011110";
        B <= "1010111010100110";
        C <= "0110001101000010";
        wait for clk_period;
        A <= "0000011100110101";
        B <= "1111010000110101";
        C <= "0000001000001000";
        wait for clk_period;
        A <= "0000111011001001";
        B <= "1100011111101000";
        C <= "1010000101101001";
        wait for clk_period;
        A <= "0011010000111010";
        B <= "1100011000011110";
        C <= "1011101000011111";
        wait for clk_period;
        A <= "1011100111010111";
        B <= "0010000011110110";
        C <= "1000000111110011";
        wait for clk_period;
        A <= "0101100110000100";
        B <= "1001001010000011";
        C <= "0101101111011111";
        wait for clk_period;
        A <= "0010001001000100";
        B <= "1110101001000100";
        C <= "1010111011111001";
        wait for clk_period;
        A <= "1111110000010100";
        B <= "0000000010011101";
        C <= "1100010011000111";
        wait for clk_period;
        A <= "1101110010001000";
        B <= "1100111011100100";
        C <= "0100100111100111";
        wait for clk_period;
        A <= "0110010100001000";
        B <= "0010101110111110";
        C <= "0111111011101111";
        wait for clk_period;
        A <= "0101101100010001";
        B <= "0000000110101001";
        C <= "0000110100000110";
        wait for clk_period;
        A <= "0001011010011110";
        B <= "0101000100101101";
        C <= "0011000001010111";
        wait for clk_period;
        A <= "0111100010110100";
        B <= "1110110101111011";
        C <= "1000010111110011";
        wait for clk_period;
        A <= "0011011001101111";
        B <= "0110011000011001";
        C <= "0010100011110010";
        wait for clk_period;
        A <= "0011101100010000";
        B <= "1111111000010010";
        C <= "1000111101100000";
        wait for clk_period;
        A <= "0000101110000011";
        B <= "1010010000111001";
        C <= "0110011011001010";
        wait for clk_period;
        A <= "1110111000010100";
        B <= "1111100011110000";
        C <= "1001011010110101";
        wait for clk_period;
        A <= "0010101111100010";
        B <= "1101010001000101";
        C <= "0000010110111011";
        wait for clk_period;
        A <= "0101101101011001";
        B <= "1110000000000110";
        C <= "1000000000011011";
        wait for clk_period;
        A <= "1101001011010110";
        B <= "1101001111011010";
        C <= "0110001111111001";
        wait for clk_period;
        A <= "0010110111111101";
        B <= "1101010011110111";
        C <= "1101110001011101";
        wait for clk_period;
        A <= "0100100011011001";
        B <= "0111000101010001";
        C <= "0010110111111010";
        wait for clk_period;
        A <= "0010011100010111";
        B <= "0001111110010011";
        C <= "1000011000110010";
        wait for clk_period;
        A <= "1111010111110100";
        B <= "1001110001111110";
        C <= "0001010100100010";
        wait for clk_period;
        A <= "0110000000010010";
        B <= "0110001001110101";
        C <= "0101011000111000";
        wait for clk_period;
        A <= "0101110000111001";
        B <= "0000111110111111";
        C <= "1101001010001011";
        wait for clk_period;
        A <= "1110111010101101";
        B <= "0001010001011001";
        C <= "0011000110110110";
        wait for clk_period;
        A <= "1101111000001100";
        B <= "0111011001100110";
        C <= "0100010110001101";
        wait for clk_period;
        A <= "0110100101110111";
        B <= "0101110101000000";
        C <= "1011110011001010";
        wait for clk_period;
        A <= "0000011010001001";
        B <= "0011001101111000";
        C <= "1110010101000011";
        wait for clk_period;
        A <= "1101001000101101";
        B <= "1000011000011110";
        C <= "0000101101001010";
        wait for clk_period;
        A <= "0000100000001000";
        B <= "1111001001010101";
        C <= "1010111010101001";
        wait for clk_period;
        A <= "0100111111011110";
        B <= "1111101011000000";
        C <= "1110100011100101";
        wait for clk_period;
        A <= "1011001100010101";
        B <= "1010110111111001";
        C <= "1001001111111000";
        wait for clk_period;
        A <= "1001101100101100";
        B <= "1101111101010011";
        C <= "0011001011110000";
        wait for clk_period;
        A <= "0110100000011010";
        B <= "1010100101101001";
        C <= "0010110111000010";
        wait for clk_period;
        A <= "1000011011000000";
        B <= "1110000000111010";
        C <= "1001100111011100";
        wait for clk_period;
        A <= "0001010011001001";
        B <= "0001000000111100";
        C <= "1001001110001110";
        wait for clk_period;
        A <= "0010100110100000";
        B <= "1010111001000010";
        C <= "1110000000100000";
        wait for clk_period;
        A <= "0110110110110011";
        B <= "0100111111111101";
        C <= "0010110110010101";
        wait for clk_period;
        A <= "1011100010000100";
        B <= "0000100100010011";
        C <= "1000110101110000";
        wait for clk_period;
        A <= "1101100110000111";
        B <= "0001101111010110";
        C <= "0001001111011111";
        wait for clk_period;
        A <= "1100001010100010";
        B <= "0110001000000001";
        C <= "0111100001110000";
        wait for clk_period;
        A <= "0000100100000101";
        B <= "0010010011100010";
        C <= "0011111100000111";
        wait for clk_period;
        A <= "0000001001001011";
        B <= "1001001111110001";
        C <= "0101010011011101";
        wait for clk_period;
        A <= "0010111001000110";
        B <= "1000001010110111";
        C <= "1010110111011001";
        wait for clk_period;
        A <= "1100111110101111";
        B <= "0110001000011101";
        C <= "1100101011110101";
        wait for clk_period;
        A <= "0011000110010111";
        B <= "0010110011100100";
        C <= "0110100001001011";
        wait for clk_period;
        A <= "1001111010000101";
        B <= "0001010101100010";
        C <= "0010000001110011";
        wait for clk_period;
        A <= "0111011001100110";
        B <= "0010100110111001";
        C <= "0011010100100111";
        wait for clk_period;
        A <= "0100011100101100";
        B <= "1101001000111011";
        C <= "0110001001111100";
        wait for clk_period;
        A <= "0101010000010110";
        B <= "0010010001011001";
        C <= "1000001111011011";
        wait for clk_period;
        A <= "1010011101000001";
        B <= "1111001011010100";
        C <= "0001010110110111";
        wait for clk_period;
        A <= "0100011101011101";
        B <= "0000010001000101";
        C <= "1110010001100100";
        wait for clk_period;
        A <= "1011110000010000";
        B <= "1101101110110110";
        C <= "0001001110001101";
        wait for clk_period;
        A <= "0010100101111101";
        B <= "0011110101010011";
        C <= "0101100100111101";
        wait for clk_period;
        A <= "0110000001011101";
        B <= "1101000110111101";
        C <= "0100011100001101";
        wait for clk_period;
        A <= "0010010011111100";
        B <= "0011011101101111";
        C <= "1101111110001111";
        wait for clk_period;
        A <= "0101010011010011";
        B <= "0010111111011100";
        C <= "0110100101010100";
        wait for clk_period;
        A <= "0110110011011001";
        B <= "1101010011000111";
        C <= "0111100011001100";
        wait for clk_period;
        A <= "0100100010101110";
        B <= "1011110001001010";
        C <= "1000110110000100";
        wait for clk_period;
        A <= "1101011111101000";
        B <= "0011010011100110";
        C <= "1101110011011101";
        wait for clk_period;
        A <= "0000000101111100";
        B <= "1010111010111101";
        C <= "0010001001011111";
        wait for clk_period;
        A <= "1101000111100010";
        B <= "0111101010000100";
        C <= "0011111110010101";
        wait for clk_period;
        A <= "0110101001000010";
        B <= "0000000110111110";
        C <= "1110000000101010";
        wait for clk_period;
        A <= "1010000010011000";
        B <= "0110010111100000";
        C <= "1110001010100011";
        wait for clk_period;
        A <= "1000100001010100";
        B <= "1100001000001010";
        C <= "1010001000010101";
        wait for clk_period;
        A <= "0011010010010000";
        B <= "1110011010000011";
        C <= "0110001000101010";
        wait for clk_period;
        A <= "1110111101110001";
        B <= "1111011111010110";
        C <= "1000110000100000";
        wait for clk_period;
        A <= "1011001110101111";
        B <= "1110100011111010";
        C <= "1000111000011101";
        wait for clk_period;
        A <= "0101100010101100";
        B <= "0101110100111111";
        C <= "0101001001101010";
        wait for clk_period;
        A <= "1000001111000011";
        B <= "1111000011100000";
        C <= "0101110111000110";
        wait for clk_period;
        A <= "1101010110101010";
        B <= "0010011011100011";
        C <= "1111000111110010";
        wait for clk_period;
        A <= "1000110101010100";
        B <= "0111111110111000";
        C <= "1101111110000111";
        wait for clk_period;
        A <= "1000011000001111";
        B <= "0100000010011011";
        C <= "0110100000000001";
        wait for clk_period;
        A <= "1001110101011111";
        B <= "0111000000010111";
        C <= "0101101110010011";
        wait for clk_period;
        A <= "0111110011010100";
        B <= "0001111110011100";
        C <= "1000110010100010";
        wait for clk_period;
        A <= "1000110110100011";
        B <= "1010101100000011";
        C <= "1011110110011010";
        wait for clk_period;
        A <= "1000011011110101";
        B <= "0110101000011011";
        C <= "0111001101010101";
        wait for clk_period;
        A <= "1100100010110111";
        B <= "0100101000101101";
        C <= "1000111000111111";
        wait for clk_period;
        A <= "1110001011100000";
        B <= "0001000000010010";
        C <= "0100101110110101";
        wait for clk_period;
        A <= "0110011001110001";
        B <= "1011000000111110";
        C <= "1110100100000101";
        wait for clk_period;
        A <= "0111001011001111";
        B <= "1110000010111101";
        C <= "0010000001111110";
        wait for clk_period;
        A <= "1010011111101110";
        B <= "1100001000110011";
        C <= "0000101011101000";
        wait for clk_period;
        A <= "0011100101010110";
        B <= "0011000011101001";
        C <= "0110101100001010";
        wait for clk_period;
        A <= "0001010110000111";
        B <= "0110010001101100";
        C <= "0001101111100000";
        wait for clk_period;
        A <= "0100011011101100";
        B <= "1111101010001010";
        C <= "0010000011111010";
        wait for clk_period;
        A <= "0111111110110111";
        B <= "0000011101000111";
        C <= "1101100111010111";
        wait for clk_period;
        A <= "0000001001011111";
        B <= "0001001100100110";
        C <= "1101010111011011";
        wait for clk_period;
        A <= "0010100110001100";
        B <= "0110010011010101";
        C <= "0011001100001110";
        wait for clk_period;
        A <= "1000110010010010";
        B <= "0010000101000001";
        C <= "1001001111011001";
        wait for clk_period;
        A <= "0011011101001000";
        B <= "0101111000100001";
        C <= "1000011011010111";
        wait for clk_period;
        A <= "0001010010000011";
        B <= "0010111110001011";
        C <= "1000101001110011";
        wait for clk_period;
        A <= "1011001011010101";
        B <= "0110111010111011";
        C <= "0101010010110010";
        wait for clk_period;
        A <= "0001101010111111";
        B <= "0101011010011101";
        C <= "0101001010001001";
        wait for clk_period;
        A <= "0100001010011101";
        B <= "0000001011000101";
        C <= "1110110111110000";
        wait for clk_period;
        A <= "1100111010000001";
        B <= "0001010001110110";
        C <= "0101010001000110";
        wait for clk_period;
        A <= "0001011001010110";
        B <= "1011111110110001";
        C <= "1001100001010100";
        wait for clk_period;
        A <= "0011111100100100";
        B <= "0001101110100101";
        C <= "1011111000100110";
        wait for clk_period;
        A <= "0010100000111010";
        B <= "1000010001000000";
        C <= "1000100100100011";
        wait for clk_period;
        A <= "0101110101000101";
        B <= "1101011101101110";
        C <= "0110000101011101";
        wait for clk_period;
        A <= "0110101111011001";
        B <= "0011011001000011";
        C <= "0001111111010111";
        wait for clk_period;
        A <= "0100100101010001";
        B <= "1110011100110110";
        C <= "1001110101111110";
        wait for clk_period;
        A <= "0011001001011000";
        B <= "1111101100101000";
        C <= "0110010000100100";
        wait for clk_period;
        A <= "0111000001100110";
        B <= "1010110011000110";
        C <= "0100001000010111";
        wait for clk_period;
        A <= "1101101111100110";
        B <= "1111111101111100";
        C <= "0001000111100111";
        wait for clk_period;
        A <= "1100101010111001";
        B <= "1001001001110110";
        C <= "1011111010111011";
        wait for clk_period;
        A <= "1010000100110000";
        B <= "1010000001100000";
        C <= "1101011101000110";
        wait for clk_period;
        A <= "1011111010001111";
        B <= "0000011100111000";
        C <= "0110101110111010";
        wait for clk_period;
        A <= "0011100111000010";
        B <= "1010101101110000";
        C <= "0111000001010011";
        wait for clk_period;
        A <= "0010101100001000";
        B <= "0010000100001100";
        C <= "0111111000011010";
        wait for clk_period;
        A <= "1111110000110011";
        B <= "0101100011101111";
        C <= "0010101011000111";
        wait for clk_period;
        A <= "1110001110101110";
        B <= "0000001010111001";
        C <= "1001100110000110";
        wait for clk_period;
        A <= "0001111000111000";
        B <= "0110001010011001";
        C <= "0110000011001111";
        wait for clk_period;
        A <= "0011001011011100";
        B <= "1100010011010001";
        C <= "1011000100001100";
        wait for clk_period;
        A <= "0111110101001000";
        B <= "1110000100001011";
        C <= "0010010011011100";
        wait for clk_period;
        A <= "0111100010101001";
        B <= "1011101111100101";
        C <= "1010111011010001";
        wait for clk_period;
        A <= "0011011110000111";
        B <= "1000011010001101";
        C <= "1111110001000010";
        wait for clk_period;
        A <= "0111001010000101";
        B <= "1100101101110010";
        C <= "1111110100110011";
        wait for clk_period;
        A <= "1111100001101001";
        B <= "0000000000100101";
        C <= "0000010101111000";
        wait for clk_period;
        A <= "0110011001110111";
        B <= "0101111111001100";
        C <= "0101110001100110";
        wait for clk_period;
        A <= "1100000000000000";
        B <= "1111010010110100";
        C <= "1100011100011100";
        wait for clk_period;
        A <= "1101111100000111";
        B <= "0000000101111011";
        C <= "0000000010001000";
        wait for clk_period;
        A <= "1001100011110000";
        B <= "0100000010000011";
        C <= "1001100111101001";
        wait for clk_period;
        A <= "0010010111101100";
        B <= "0101000001110000";
        C <= "1000000110111110";
        wait for clk_period;
        A <= "1011011111100001";
        B <= "1011000111110001";
        C <= "0100100100100000";
        wait for clk_period;
        A <= "1101001000110010";
        B <= "1100100111011101";
        C <= "0011111000010101";
        wait for clk_period;
        A <= "1100110100011001";
        B <= "0011101111001010";
        C <= "0101000110111010";
        wait for clk_period;
        A <= "1011101011000110";
        B <= "1011101111111001";
        C <= "0000100111000111";
        wait for clk_period;
        A <= "1001110100111000";
        B <= "1110011000110010";
        C <= "1000001000000101";
        wait for clk_period;
        A <= "0110100001000100";
        B <= "1011000000111101";
        C <= "0100010000100101";
        wait for clk_period;
        A <= "0011011101101111";
        B <= "1100011111101100";
        C <= "1100001001110110";
        wait for clk_period;
        A <= "1001011000111100";
        B <= "0000011010000101";
        C <= "1000100110110010";
        wait for clk_period;
        A <= "1111001101001011";
        B <= "0011110010010101";
        C <= "1001010000011101";
        wait for clk_period;
        A <= "0010110001110110";
        B <= "0100001001101110";
        C <= "0110101111101010";
        wait for clk_period;
        A <= "0010011001011110";
        B <= "1101000101110101";
        C <= "0111011100001001";
        wait for clk_period;
        A <= "1010100101101011";
        B <= "0100010000000111";
        C <= "0101010000000100";
        wait for clk_period;
        A <= "0111010011001001";
        B <= "0010011100100111";
        C <= "1101100001001110";
        wait for clk_period;
        A <= "1111000000001111";
        B <= "1011110001100101";
        C <= "0001100000110000";
        wait for clk_period;
        A <= "0110111110011001";
        B <= "0101111111101100";
        C <= "1100110011110000";
        wait for clk_period;
        A <= "1010001011010100";
        B <= "1111110011001010";
        C <= "1101111100010111";
        wait for clk_period;
        A <= "0101001001011001";
        B <= "1011010110010100";
        C <= "0111010111101111";
        wait for clk_period;
        A <= "0110000001011011";
        B <= "1101100011011010";
        C <= "1000001001001000";
        wait for clk_period;
        A <= "1001001100011000";
        B <= "0011110111110101";
        C <= "1100001111111010";
        wait for clk_period;
        A <= "0111000011110010";
        B <= "1111000100111110";
        C <= "0111001001101010";
        wait for clk_period;
        A <= "0100010010100010";
        B <= "1010101101010101";
        C <= "1111111110010101";
        wait for clk_period;
        A <= "1100110100111111";
        B <= "0000110111000011";
        C <= "1010101001111111";
        wait for clk_period;
        A <= "1101000101010011";
        B <= "1111000010011011";
        C <= "0100110101010111";
        wait for clk_period;
        A <= "1011100000010000";
        B <= "0101101110100000";
        C <= "0100100000010000";
        wait for clk_period;
        A <= "1111011010000010";
        B <= "0101111001101001";
        C <= "0101000001110110";
        wait for clk_period;
        A <= "1101000010000111";
        B <= "0100101011000100";
        C <= "1011110000110010";
        wait for clk_period;
        A <= "0001010101001100";
        B <= "0001110110100100";
        C <= "0111010000000011";
        wait for clk_period;
        A <= "1101011000001001";
        B <= "0110001010101010";
        C <= "0011110100011010";
        wait for clk_period;
        A <= "1100111000000111";
        B <= "1110110110101011";
        C <= "1011000101100001";
        wait for clk_period;
        A <= "0010101001011001";
        B <= "0101101000111101";
        C <= "1010110001000001";
        wait for clk_period;
        A <= "0011111000000101";
        B <= "0111100010011100";
        C <= "0000110011011101";
        wait for clk_period;
        A <= "0011110110111101";
        B <= "0111011001100110";
        C <= "0001001001011101";
        wait for clk_period;
        A <= "1110100100101100";
        B <= "0110101101001110";
        C <= "0101000100101101";
        wait for clk_period;
        A <= "1001100001110001";
        B <= "0011010111110110";
        C <= "0111100010110110";
        wait for clk_period;
        A <= "1000001110101110";
        B <= "1001000010110101";
        C <= "1010001001100101";
        wait for clk_period;
        A <= "1010110111111110";
        B <= "0011110100101001";
        C <= "0010100000101000";
        wait for clk_period;
        A <= "1010100000010010";
        B <= "1101100000111000";
        C <= "0100101100001101";
        wait for clk_period;
        A <= "1101001110110111";
        B <= "1100100001000010";
        C <= "0101100101010010";
        wait for clk_period;
        A <= "0000101101000110";
        B <= "1010010000101110";
        C <= "0011100010111010";
        wait for clk_period;
        A <= "0010101101000100";
        B <= "1001001100100001";
        C <= "0001010001100011";
        wait for clk_period;
        A <= "1110010000111100";
        B <= "1001011110000101";
        C <= "0110111101100011";
        wait for clk_period;
        A <= "0101100001001000";
        B <= "0110111100000110";
        C <= "0011001100001101";
        wait for clk_period;
        A <= "1011111110001110";
        B <= "0101010100010000";
        C <= "1110100011101111";
        wait for clk_period;
        A <= "1010000110111000";
        B <= "0010101100101101";
        C <= "1111011111000110";
        wait for clk_period;
        A <= "1110100010111100";
        B <= "0110010000011001";
        C <= "1011100100011111";
        wait for clk_period;
        A <= "0111001101100101";
        B <= "1101010100011001";
        C <= "0100010010000001";
        wait for clk_period;
        A <= "0100111111011111";
        B <= "1001110001011111";
        C <= "0011110000011101";
        wait for clk_period;
        A <= "1100110111110101";
        B <= "1010000100100110";
        C <= "1101110001001111";
        wait for clk_period;
        A <= "0001001011101101";
        B <= "1110100000000110";
        C <= "0111101011010000";
        wait for clk_period;
        A <= "1001000111011111";
        B <= "1111111100101011";
        C <= "0111101110000100";
        wait for clk_period;
        A <= "1101001100101000";
        B <= "0011000001001111";
        C <= "1110001011100000";
        wait for clk_period;
        A <= "1111110011100111";
        B <= "1110111110001011";
        C <= "1100001011100111";
        wait for clk_period;
        A <= "0000110110010010";
        B <= "0001011110110000";
        C <= "1110011000011101";
        wait for clk_period;
        A <= "0110001110001001";
        B <= "0110111100101111";
        C <= "1011001000100100";
        wait for clk_period;
        A <= "1000011101101110";
        B <= "1011001101110111";
        C <= "0110100010001111";
        wait for clk_period;
        A <= "0001111000101111";
        B <= "1110100100001100";
        C <= "0000110011000101";
        wait for clk_period;
        A <= "0100011010011101";
        B <= "1001010100011001";
        C <= "0010101011001111";
        wait for clk_period;
        A <= "1001101111100001";
        B <= "1110010100110110";
        C <= "1101000000010011";
        wait for clk_period;
        A <= "1010110100000010";
        B <= "1010110111011110";
        C <= "1011111011000101";
        wait for clk_period;
        A <= "0110100010000111";
        B <= "0000010101101111";
        C <= "1110110001011000";
        wait for clk_period;
        A <= "1110111100011001";
        B <= "0000100101000000";
        C <= "1001000010101011";
        wait for clk_period;
        A <= "1101010010111101";
        B <= "0100101110000101";
        C <= "0110110000001011";
        wait for clk_period;
        A <= "1011101100011011";
        B <= "1111110011100100";
        C <= "0011101101000110";
        wait for clk_period;
        A <= "1101010110001110";
        B <= "1001001101001001";
        C <= "0001010001011101";
        wait for clk_period;
        A <= "1011111111011000";
        B <= "0100011111100100";
        C <= "0011100000000101";
        wait for clk_period;
        A <= "1001011001001110";
        B <= "1110000100101110";
        C <= "1110011001110011";
        wait for clk_period;
        A <= "1110110100111001";
        B <= "0100100111100011";
        C <= "1011110010101000";
        wait for clk_period;
        A <= "0000000011110101";
        B <= "0011000011101011";
        C <= "0110011001010111";
        wait for clk_period;
        A <= "0101000101100010";
        B <= "0011101000100100";
        C <= "0000101101111000";
        wait for clk_period;
        A <= "0100000001101110";
        B <= "1010001001110001";
        C <= "0010111011100001";
        wait for clk_period;
        A <= "1111010010010011";
        B <= "0100001100000111";
        C <= "0110001010100011";
        wait for clk_period;
        A <= "1101001100100000";
        B <= "1010010111011000";
        C <= "1010010111111010";
        wait for clk_period;
        A <= "0001001111101111";
        B <= "1000001100011011";
        C <= "0100010010001101";
        wait for clk_period;
        A <= "1101011110101111";
        B <= "0100001110101100";
        C <= "1011111111111111";
        wait for clk_period;
        A <= "1111101010111010";
        B <= "1111110111010001";
        C <= "0111000001001010";
        wait for clk_period;
        A <= "1001001010110000";
        B <= "0010101010100101";
        C <= "1011111101010110";
        wait for clk_period;
        A <= "0011100010011001";
        B <= "0110010101101010";
        C <= "0001110001101000";
        wait for clk_period;
        A <= "1011000010110001";
        B <= "1100111100010001";
        C <= "0000001001101011";
        wait for clk_period;
        A <= "1100100111101110";
        B <= "0011001110110100";
        C <= "1011100100100110";
        wait for clk_period;
        A <= "1011010001011110";
        B <= "0010001011111011";
        C <= "1010001111010111";
        wait for clk_period;
        A <= "1011110110101000";
        B <= "1010011110011001";
        C <= "0110101101101110";
        wait for clk_period;
        A <= "1011010111000101";
        B <= "1111011111101100";
        C <= "1110011001010101";
        wait for clk_period;
        A <= "1100100110010010";
        B <= "0111001111010101";
        C <= "1111000011010100";
        wait for clk_period;
        A <= "1111100000110101";
        B <= "0101101110110011";
        C <= "1001000101111110";
        wait for clk_period;
        A <= "1011001110010001";
        B <= "1111010100100000";
        C <= "1101110110101001";
        wait for clk_period;
        A <= "1000011111100111";
        B <= "0001001100000001";
        C <= "1011011001000110";
        wait for clk_period;
        A <= "0101011101011010";
        B <= "0110100101000101";
        C <= "1001111101000000";
        wait for clk_period;
        A <= "0011000111111101";
        B <= "0011010010111000";
        C <= "1100101001010101";
        wait for clk_period;
        A <= "1100001101110110";
        B <= "0111010101101100";
        C <= "0000001110010011";
        wait for clk_period;
        A <= "0110100110001011";
        B <= "1110111111010010";
        C <= "1001110000100000";
        wait for clk_period;
        A <= "1011000000011111";
        B <= "1101011000110100";
        C <= "0110010100010111";
        wait for clk_period;
        A <= "0011011000000010";
        B <= "1011011001111100";
        C <= "1101110011001101";
        wait for clk_period;
        A <= "1010100011101101";
        B <= "0010011100111101";
        C <= "1001000010111001";
        wait for clk_period;
        A <= "0111111001101000";
        B <= "0101011011000111";
        C <= "1000110100110101";
        wait for clk_period;
        A <= "0000111101010100";
        B <= "0010011011111110";
        C <= "0100110101011100";
        wait for clk_period;
        A <= "1111000011011100";
        B <= "0001001110100010";
        C <= "1000000010011110";
        wait for clk_period;
        A <= "1010000001111010";
        B <= "1001110111110011";
        C <= "0111110101110000";
        wait for clk_period;
        A <= "1011001000000010";
        B <= "0001100001101001";
        C <= "1110101100111010";
        wait for clk_period;
        A <= "1011010101111110";
        B <= "0100010011000001";
        C <= "0101101001000110";
        wait for clk_period;
        A <= "1100101001110111";
        B <= "1110100110010100";
        C <= "1001000101111101";
        wait for clk_period;
        A <= "1011010000110101";
        B <= "0100001010000010";
        C <= "1001000011100111";
        wait for clk_period;
        A <= "1101011111111101";
        B <= "1011100101001001";
        C <= "0111110010001100";
        wait for clk_period;
        A <= "1000000111011100";
        B <= "1100000100010101";
        C <= "0101111010111000";
        wait for clk_period;
        A <= "0101001000000000";
        B <= "0000010111011100";
        C <= "1010111111000000";
        wait for clk_period;
        A <= "1101011001101100";
        B <= "0011011101010011";
        C <= "1000011001010000";
        wait for clk_period;
        A <= "1111110100101000";
        B <= "0110011010100110";
        C <= "1010001010101001";
        wait for clk_period;
        A <= "0001101101100000";
        B <= "1110100100100010";
        C <= "0111000011000000";
        wait for clk_period;
        A <= "0111101010001001";
        B <= "0101011001001011";
        C <= "1110011111111001";
        wait for clk_period;
        A <= "0001010000100111";
        B <= "1001010011010100";
        C <= "0011111111000111";
        wait for clk_period;
        A <= "0011111111010101";
        B <= "0110110000010111";
        C <= "1110001010101110";
        wait for clk_period;
        A <= "0010111010011110";
        B <= "0011111011100010";
        C <= "0010010010000001";
        wait for clk_period;
        A <= "0110111000101110";
        B <= "0111100001100011";
        C <= "0100111010010100";
        wait for clk_period;
        A <= "0100101101011000";
        B <= "0101000111001111";
        C <= "1100101101110011";
        wait for clk_period;
        A <= "1011110000110000";
        B <= "1101100110100100";
        C <= "0000010100000000";
        wait for clk_period;
        A <= "1100000111010011";
        B <= "0000010111110001";
        C <= "1010000100101100";
        wait for clk_period;
        A <= "1001001000100000";
        B <= "0110011001000100";
        C <= "1110011011100000";
        wait for clk_period;
        A <= "1010111101011101";
        B <= "0101011011100010";
        C <= "0101111000100100";
        wait for clk_period;
        A <= "0010011101010100";
        B <= "0001100011001101";
        C <= "1110101100010100";
        wait for clk_period;
        A <= "0001110011000001";
        B <= "0010111001100010";
        C <= "1001010001001101";
        wait for clk_period;
        A <= "1100101111001111";
        B <= "1010011010111111";
        C <= "0100111010010001";
        wait for clk_period;
        A <= "0101000011101111";
        B <= "0100001001010010";
        C <= "1111000101101011";
        wait for clk_period;
        A <= "1100101101111010";
        B <= "0100111010111100";
        C <= "0101101101110111";
        wait for clk_period;
        A <= "1001000000100111";
        B <= "1001100000001010";
        C <= "0100000000010011";
        wait for clk_period;
        A <= "0000110001100000";
        B <= "1001010101110101";
        C <= "0100000110101100";
        wait for clk_period;
        A <= "1100010000101111";
        B <= "1111100101011110";
        C <= "0001000001000110";
        wait for clk_period;
        A <= "0001100111000111";
        B <= "1110101111000110";
        C <= "0001011111001101";
        wait for clk_period;
        A <= "0000011101111011";
        B <= "1010001100011101";
        C <= "0111011001011111";
        wait for clk_period;
        A <= "1000011100000011";
        B <= "0001000011001001";
        C <= "1101001001000100";
        wait for clk_period;
        A <= "0000000010110110";
        B <= "1010101010011100";
        C <= "0111000011000010";
        wait for clk_period;
        A <= "1100000011000011";
        B <= "0101001000011110";
        C <= "1100001110110000";
        wait for clk_period;
        A <= "0101000110111101";
        B <= "0011000101010111";
        C <= "0111011000011010";
        wait for clk_period;
        A <= "0110110100010001";
        B <= "1000101100010101";
        C <= "1011100101011111";
        wait for clk_period;
        A <= "1100010100101000";
        B <= "0101011000001011";
        C <= "1100111101001011";
        wait for clk_period;
        A <= "1111110111101011";
        B <= "1101111010111011";
        C <= "0000101111100011";
        wait for clk_period;
        A <= "0001010101011111";
        B <= "0111001000000101";
        C <= "1010110100001101";
        wait for clk_period;
        A <= "0011101000011011";
        B <= "1111001010011111";
        C <= "0011110011111101";
        wait for clk_period;
        A <= "0000001101110111";
        B <= "1101110101100111";
        C <= "1010101110010101";
        wait for clk_period;
        A <= "1011110010010100";
        B <= "0101001100001100";
        C <= "1100011111100001";
        wait for clk_period;
        A <= "1001011100100100";
        B <= "0011100011100010";
        C <= "1101011111000110";
        wait for clk_period;
        A <= "0100001011010110";
        B <= "1100010000101001";
        C <= "1100011010011011";
        wait for clk_period;
        A <= "0110110111011100";
        B <= "1011011110001001";
        C <= "1111000011011011";
        wait for clk_period;
        A <= "0001111011101111";
        B <= "0110010001101001";
        C <= "1101010110110000";
        wait for clk_period;
        A <= "0000101011110010";
        B <= "0000010100011010";
        C <= "0110000000110110";
        wait for clk_period;
        A <= "0101110001010110";
        B <= "0010010011000010";
        C <= "1101000100110011";
        wait for clk_period;
        A <= "1011101011011010";
        B <= "0101011100101101";
        C <= "0101100111011010";
        wait for clk_period;
        A <= "1000100111100010";
        B <= "1101110011111110";
        C <= "1111111000001100";
        wait for clk_period;
        A <= "0100001101011011";
        B <= "1101110010110110";
        C <= "1100110110010010";
        wait for clk_period;
        A <= "0011000101111011";
        B <= "1000110100011010";
        C <= "1111001110011000";
        wait for clk_period;
        A <= "0101100101010000";
        B <= "0011100101100111";
        C <= "1001010011010000";
        wait for clk_period;
        A <= "0100000010111011";
        B <= "1000001011101000";
        C <= "1101110100111111";
        wait for clk_period;
        A <= "1001111001100010";
        B <= "1101000011001010";
        C <= "1101011010011000";
        wait for clk_period;
        A <= "1010000100011100";
        B <= "1111000011001010";
        C <= "0111100111001001";
        wait for clk_period;
        A <= "1110101110110011";
        B <= "1111000000000110";
        C <= "0110011011001010";
        wait for clk_period;
        A <= "1001000000000011";
        B <= "0101001100100010";
        C <= "0110010011001011";
        wait for clk_period;
        A <= "0100011101100101";
        B <= "1110100010110110";
        C <= "1001100000110001";
        wait for clk_period;
        A <= "1010110000101101";
        B <= "1110000000001110";
        C <= "0011111010001110";
        wait for clk_period;
        A <= "0111101011111000";
        B <= "0100111100001101";
        C <= "0010111111001011";
        wait for clk_period;
        A <= "1010101010010101";
        B <= "1110111111110101";
        C <= "1001101100000110";
        wait for clk_period;
        A <= "0111101010100001";
        B <= "1001101101010101";
        C <= "1000100010101111";
        wait for clk_period;
        A <= "1110100110101101";
        B <= "0101011010101000";
        C <= "1011000101011100";
        wait for clk_period;
        A <= "1010111001011110";
        B <= "0010010010100111";
        C <= "1011011100100101";
        wait for clk_period;
        A <= "1101110001111001";
        B <= "1110001010110100";
        C <= "0110010000011011";
        wait for clk_period;
        A <= "1101010100010011";
        B <= "1010000001101000";
        C <= "0000110101101100";
        wait for clk_period;
        A <= "1111000000011000";
        B <= "1101011011111101";
        C <= "1101001110001010";
        wait for clk_period;
        A <= "0001000100010000";
        B <= "1011111110001010";
        C <= "0111110010001100";
        wait for clk_period;
        A <= "0011100000010001";
        B <= "1010000101010001";
        C <= "1101010010011100";
        wait for clk_period;
        A <= "0011101111101101";
        B <= "0111001101111100";
        C <= "0010011101100011";
        wait for clk_period;
        A <= "1010100010011010";
        B <= "0011110001010111";
        C <= "1101011000001000";
        wait for clk_period;
        A <= "1110011001010101";
        B <= "1010100011101100";
        C <= "1110101111100000";
        wait for clk_period;
        A <= "0110000000001011";
        B <= "1110010100101001";
        C <= "0010001011011010";
        wait for clk_period;
        A <= "0100111001000111";
        B <= "1001001111101001";
        C <= "0100111101010001";
        wait for clk_period;
        A <= "0111010011111111";
        B <= "1101101011101111";
        C <= "1000011011000010";
        wait for clk_period;
        A <= "0010110101001111";
        B <= "1100110110011110";
        C <= "0111010100110110";
        wait for clk_period;
        A <= "1010000110100111";
        B <= "1100101101010011";
        C <= "0100001010110100";
        wait for clk_period;
        A <= "0010011100000111";
        B <= "0100101001111111";
        C <= "1110100100000010";
        wait for clk_period;
        A <= "1011100000001001";
        B <= "1010011000000101";
        C <= "1010111001101001";
        wait for clk_period;
        A <= "1110010000111101";
        B <= "0100101011110111";
        C <= "0100101000100001";
        wait for clk_period;
        A <= "1100010110100110";
        B <= "1000111100101111";
        C <= "0010000100011000";
        wait for clk_period;
        A <= "1111111100111000";
        B <= "0011000111001110";
        C <= "0100001010010100";
        wait for clk_period;
        A <= "0110010111000100";
        B <= "0101011100010100";
        C <= "0000110100101110";
        wait for clk_period;
        A <= "0100100111011010";
        B <= "1000110000000101";
        C <= "1100011101111010";
        wait for clk_period;
        A <= "1101101010010100";
        B <= "0001001000111010";
        C <= "0110100100001101";
        wait for clk_period;
        A <= "0001100000000011";
        B <= "1001000100101011";
        C <= "0110110101100101";
        wait for clk_period;
        A <= "1101011010011111";
        B <= "1110110001100000";
        C <= "1111101010001101";
        wait for clk_period;
        A <= "0011000111010001";
        B <= "1101110000010110";
        C <= "0011101111001011";
        wait for clk_period;
        A <= "0001100000010010";
        B <= "1110111110010101";
        C <= "1110000001011111";
        wait for clk_period;
        A <= "0100111110001011";
        B <= "0100001101011000";
        C <= "0111110110110000";
        wait for clk_period;
        A <= "0000010011011001";
        B <= "1100001111111111";
        C <= "1100111000001100";
        wait for clk_period;
        A <= "0000011011000001";
        B <= "1011101100011000";
        C <= "1000010001011011";
        wait for clk_period;
        A <= "0100011100000011";
        B <= "1100011000100011";
        C <= "1001100100101010";
        wait for clk_period;
        A <= "0111101011000110";
        B <= "0100101011010101";
        C <= "1100001101011100";
        wait for clk_period;
        A <= "0001000111100011";
        B <= "0110101001000101";
        C <= "0111001010010010";
        wait for clk_period;
        A <= "1110101100111100";
        B <= "0100101010000111";
        C <= "1000110101000000";
        wait for clk_period;
        A <= "1110100000000100";
        B <= "0100100011111111";
        C <= "1101100111110001";
        wait for clk_period;
        A <= "0010011111100000";
        B <= "0111110111111100";
        C <= "1010000100101100";
        wait for clk_period;
        A <= "0100001110111110";
        B <= "1100101001111000";
        C <= "1111011100010111";
        wait for clk_period;
        A <= "1001111100101100";
        B <= "0111001110101101";
        C <= "1111110111010101";
        wait for clk_period;
        A <= "0011111101001000";
        B <= "0010101011110001";
        C <= "1011010000011001";
        wait for clk_period;
        A <= "0000111000100000";
        B <= "0001000100011010";
        C <= "0000001101111101";
        wait for clk_period;
        A <= "1000010111100100";
        B <= "1011101011001111";
        C <= "0110011100010101";
        wait for clk_period;
        A <= "1010001011000011";
        B <= "1100001010101100";
        C <= "0011100010000110";
        wait for clk_period;
        A <= "0000100101110010";
        B <= "1110000110110111";
        C <= "0010101000110011";
        wait for clk_period;
        A <= "1010111101001010";
        B <= "1110001101100100";
        C <= "0110000110010011";
        wait for clk_period;
        A <= "1001101001010100";
        B <= "0110011000011001";
        C <= "0000000110101111";
        wait for clk_period;
        A <= "0001100000101010";
        B <= "0110111111100101";
        C <= "0101001000101010";
        wait for clk_period;
        A <= "0001000101000011";
        B <= "0000110110110000";
        C <= "0010001001110001";
        wait for clk_period;
        A <= "1010110110000101";
        B <= "0101011010000101";
        C <= "0000101000101011";
        wait for clk_period;
        A <= "0011111011001011";
        B <= "1000100001110010";
        C <= "1000010101100011";
        wait for clk_period;
        A <= "1111101000101110";
        B <= "1001000101001011";
        C <= "0100000000100101";
        wait for clk_period;
        A <= "0110000111010110";
        B <= "1001100111001000";
        C <= "1110101100001110";
        wait for clk_period;
        A <= "1101010101111010";
        B <= "0100101110010100";
        C <= "0010100100011111";
        wait for clk_period;
        A <= "0011100110100011";
        B <= "0011100110101110";
        C <= "1010111000011001";
        wait for clk_period;
        A <= "1001000000010010";
        B <= "1001110101010111";
        C <= "1111001001100011";
        wait for clk_period;
        A <= "0000000111110010";
        B <= "0101111110110101";
        C <= "1111111000101100";
        wait for clk_period;
        A <= "0101000101011001";
        B <= "1011001011000110";
        C <= "0100100000010110";
        wait for clk_period;
        A <= "1011101000000110";
        B <= "0011100011000000";
        C <= "0100110011110100";
        wait for clk_period;
        A <= "1110110111101001";
        B <= "1001010010001110";
        C <= "0001100100110000";
        wait for clk_period;
        A <= "0100000011100101";
        B <= "1010001100110010";
        C <= "1101011101011101";
        wait for clk_period;
        A <= "1111010100100000";
        B <= "0011001100010011";
        C <= "1110000100111100";
        wait for clk_period;
        A <= "1100101001111011";
        B <= "1001101000001101";
        C <= "0011010001100010";
        wait for clk_period;
        A <= "1100101000011101";
        B <= "0110011010111011";
        C <= "0101011100011111";
        wait for clk_period;
        A <= "1000111110110000";
        B <= "1011011000000111";
        C <= "1010110001100011";
        wait for clk_period;
        A <= "1100101000100111";
        B <= "1001101111010010";
        C <= "1010010011101011";
        wait for clk_period;
        A <= "0110111000111110";
        B <= "1011110100000100";
        C <= "0100111100110110";
        wait for clk_period;
        A <= "0100011000011111";
        B <= "1101100000100000";
        C <= "0001100000110001";
        wait for clk_period;
        A <= "1010011001100000";
        B <= "0000101111010101";
        C <= "1011101101000111";
        wait for clk_period;
        A <= "0000001001000101";
        B <= "0000100011100011";
        C <= "0100101100000000";
        wait for clk_period;
        A <= "1100101110101001";
        B <= "1000010101000001";
        C <= "0100101100010101";
        wait for clk_period;
        A <= "1001111110010011";
        B <= "1110000001011001";
        C <= "1011000100011000";
        wait for clk_period;
        A <= "0100011001100111";
        B <= "0100010110011001";
        C <= "1011000001100101";
        wait for clk_period;
        A <= "1100001000000010";
        B <= "0110100000100000";
        C <= "1011101110100011";
        wait for clk_period;
        A <= "0100101111010001";
        B <= "0000101111000000";
        C <= "1110000111000111";
        wait for clk_period;
        A <= "1000110001010111";
        B <= "1010011001000010";
        C <= "0111101001101101";
        wait for clk_period;
        A <= "1110011000001011";
        B <= "0011000111001000";
        C <= "1011111111000001";
        wait for clk_period;
        A <= "1111000110000001";
        B <= "0110000010101010";
        C <= "0011111100000011";
        wait for clk_period;
        A <= "1110110001110000";
        B <= "0110010010110010";
        C <= "1110111001110101";
        wait for clk_period;
        A <= "0100110010000000";
        B <= "0101001101000010";
        C <= "1001000010001111";
        wait for clk_period;
        A <= "0110100101010100";
        B <= "0110110101011011";
        C <= "0000101110110011";
        wait for clk_period;
        A <= "1000000011001001";
        B <= "1110100000111100";
        C <= "0100111100000011";
        wait for clk_period;
        A <= "1011101100100101";
        B <= "1011000010111111";
        C <= "0010000001111100";
        wait for clk_period;
        A <= "0011011010010110";
        B <= "1000011111110111";
        C <= "1111001111101000";
        wait for clk_period;
        A <= "1000011000100110";
        B <= "1000000000010011";
        C <= "1110101010100011";
        wait for clk_period;
        A <= "0000100010000000";
        B <= "0111100110100000";
        C <= "0010010101101011";
        wait for clk_period;
        A <= "1101100110101110";
        B <= "0011001101101101";
        C <= "1100110110011011";
        wait for clk_period;
        A <= "1010111010000011";
        B <= "1111100111101011";
        C <= "1101110011101100";
        wait for clk_period;
        A <= "0111001000011000";
        B <= "0000011101010011";
        C <= "1000010000111101";
        wait for clk_period;
        A <= "0100100101111101";
        B <= "1001110010111100";
        C <= "0100000111110101";
        wait for clk_period;
        A <= "1111000000010111";
        B <= "0110000000101000";
        C <= "0001111000110001";
        wait for clk_period;
        A <= "0101110000001111";
        B <= "1111110110010100";
        C <= "1010000100010001";
        wait for clk_period;
        A <= "1100100000000010";
        B <= "1000100010100111";
        C <= "0000101001001011";
        wait for clk_period;
        A <= "1010000101011010";
        B <= "1111011010101111";
        C <= "0000100111101001";
        wait for clk_period;
        A <= "0001000100000100";
        B <= "0011011010010101";
        C <= "1000001010011010";
        wait for clk_period;
        A <= "0001100101010111";
        B <= "1101100010000110";
        C <= "0101000011100100";
        wait for clk_period;
        A <= "1100101111011100";
        B <= "1000010010000110";
        C <= "0111110000001100";
        wait for clk_period;
        A <= "0101101011001011";
        B <= "0011011011100001";
        C <= "1010101101100110";
        wait for clk_period;
        A <= "0010100010101001";
        B <= "1110110010001110";
        C <= "1010110011111000";
        wait for clk_period;
        A <= "1001011011110000";
        B <= "1110000100011000";
        C <= "1001101001011101";
        wait for clk_period;
        A <= "1110100001000011";
        B <= "1000011001111011";
        C <= "1110111000100100";
        wait for clk_period;
        A <= "0000010001000011";
        B <= "0000101011101010";
        C <= "1111101100011001";
        wait for clk_period;
        A <= "0111000100000110";
        B <= "1011111101101000";
        C <= "0101011010010011";
        wait for clk_period;
        A <= "0001000011001101";
        B <= "0001101011100101";
        C <= "1110100011111001";
        wait for clk_period;
        A <= "0101011101000001";
        B <= "1000101110101100";
        C <= "0011111000011011";
        wait for clk_period;
        A <= "0100001010001100";
        B <= "0001011011110010";
        C <= "1101111000000111";
        wait for clk_period;
        A <= "0001011111100100";
        B <= "1001011000110010";
        C <= "0001001000001111";
        wait for clk_period;
        A <= "0010110110100100";
        B <= "1100111000110011";
        C <= "0110000001100001";
        wait for clk_period;
        A <= "0100010001101001";
        B <= "1001000000000101";
        C <= "1000100011001100";
        wait for clk_period;
        A <= "1000000101100010";
        B <= "0110010010111001";
        C <= "1001000001001100";
        wait for clk_period;
        A <= "1000010110110010";
        B <= "0110110101001000";
        C <= "0100010101100100";
        wait for clk_period;
        A <= "0101001010010111";
        B <= "0011100101110010";
        C <= "0000101111101010";
        wait for clk_period;
        A <= "0110110110101001";
        B <= "0100010000010000";
        C <= "1001011101110101";
        wait for clk_period;
        A <= "1001110100011000";
        B <= "1011101000100001";
        C <= "0101110111110100";
        wait for clk_period;
        A <= "1101111111111100";
        B <= "0110000100101010";
        C <= "0100001010111010";
        wait for clk_period;
        A <= "0101011000111101";
        B <= "1111111001010101";
        C <= "1100001011101110";
        wait for clk_period;
        A <= "1111000111001000";
        B <= "0010010011111100";
        C <= "0001110010101011";
        wait for clk_period;
        A <= "0010011010011001";
        B <= "1010100000011010";
        C <= "1110101110101111";
        wait for clk_period;
        A <= "0000001011000100";
        B <= "0111111000111001";
        C <= "0110010100111100";
        wait for clk_period;
        A <= "0011100011011110";
        B <= "0110111010110111";
        C <= "0100011000101101";
        wait for clk_period;
        A <= "1111011001000111";
        B <= "0100001100001110";
        C <= "0110000110101000";
        wait for clk_period;
        A <= "0100011011011110";
        B <= "0001000110001101";
        C <= "1100100111101111";
        wait for clk_period;
        A <= "1000001111001000";
        B <= "1000000110000000";
        C <= "1100001100000000";
        wait for clk_period;
        A <= "1001110110100110";
        B <= "0000110000010101";
        C <= "0000001101100001";
        wait for clk_period;
        A <= "1111011110010011";
        B <= "1111100010011000";
        C <= "0000100111111010";
        wait for clk_period;
        A <= "0001101011101111";
        B <= "0110100000100001";
        C <= "0110011100000110";
        wait for clk_period;
        A <= "0010101111110000";
        B <= "0111100100011001";
        C <= "0101010001000010";
        wait for clk_period;
        A <= "1110111011111011";
        B <= "1001101111111010";
        C <= "1001110000111010";
        wait for clk_period;
        A <= "1000110011011010";
        B <= "1010101001100000";
        C <= "0001010100111000";
        wait for clk_period;
        A <= "0011100101001100";
        B <= "0010011100111000";
        C <= "0101001100101011";
        wait for clk_period;
        A <= "0011100100011010";
        B <= "0011101111001001";
        C <= "0100001010101100";
        wait for clk_period;
        A <= "1100011000100001";
        B <= "0010100000001000";
        C <= "1010111010001010";
        wait for clk_period;
        A <= "0000111000101111";
        B <= "1100101110001110";
        C <= "0001000000110111";
        wait for clk_period;
        A <= "1000001011110110";
        B <= "0110101100000101";
        C <= "0110000000011011";
        wait for clk_period;
        A <= "0010011010100100";
        B <= "0111010101011100";
        C <= "0100010110111100";
        wait for clk_period;
        A <= "1011111001111001";
        B <= "1001110000101110";
        C <= "0001000000010111";
        wait for clk_period;
        A <= "1111011001011110";
        B <= "0110110110011100";
        C <= "1100011000011000";
        wait for clk_period;
        A <= "1101010010111000";
        B <= "1010001001111111";
        C <= "1101101111001011";
        wait for clk_period;
        A <= "0000011110000000";
        B <= "0000000010100111";
        C <= "1101111111000110";
        wait for clk_period;
        A <= "1100001111011011";
        B <= "1111110101001101";
        C <= "1011101101100111";
        wait for clk_period;
        A <= "0011111101100100";
        B <= "0100100011001011";
        C <= "0101111010111100";
        wait for clk_period;
        A <= "1111001110000111";
        B <= "0100100010101011";
        C <= "1000100000001001";
        wait for clk_period;
        A <= "0001101101100110";
        B <= "0001101000010100";
        C <= "0101101110010100";
        wait for clk_period;
        A <= "0011101011011000";
        B <= "1101001110010010";
        C <= "1111001110110110";
        wait for clk_period;
        A <= "1010010001010010";
        B <= "0010111010100110";
        C <= "1100000110110100";
        wait for clk_period;
        A <= "1011001000001010";
        B <= "1000100111110111";
        C <= "1000111010000100";
        wait for clk_period;
        A <= "1001001010100010";
        B <= "0010100010001000";
        C <= "0110001110011010";
        wait for clk_period;
        A <= "0111110000111001";
        B <= "0010010100111110";
        C <= "1011110010001111";
        wait for clk_period;
        A <= "0110100100111110";
        B <= "0011110111110111";
        C <= "1010111100001010";
        wait for clk_period;
        A <= "1000001111101111";
        B <= "1111011000000100";
        C <= "1110100100101110";
        wait for clk_period;
        A <= "1011101001010001";
        B <= "1011111000101111";
        C <= "1111111010101111";
        wait for clk_period;
        A <= "1100110111111100";
        B <= "1100001000001101";
        C <= "0100000010001101";
        wait for clk_period;
        A <= "0000110110010100";
        B <= "0111001011100111";
        C <= "1010111111010001";
        wait for clk_period;
        A <= "0101001011110100";
        B <= "1011100011010110";
        C <= "1010011110010000";
        wait for clk_period;
        A <= "0100110001110010";
        B <= "0101010100000011";
        C <= "1011011100010100";
        wait for clk_period;
        A <= "0101000110101001";
        B <= "0011111000110010";
        C <= "0110010101011011";
        wait for clk_period;
        A <= "1110010110100100";
        B <= "0001001101000000";
        C <= "1011100011011100";
        wait for clk_period;
        A <= "0000110100101001";
        B <= "1011101101111000";
        C <= "0011000001011100";
        wait for clk_period;
        A <= "1110110011111110";
        B <= "0101100000100001";
        C <= "1110110101100001";
        wait for clk_period;
        A <= "1000100011000010";
        B <= "0110110111001010";
        C <= "1100111001010111";
        wait for clk_period;
        A <= "0011100111100011";
        B <= "1111000111000101";
        C <= "0110011000100011";
        wait for clk_period;
        A <= "0011000011100100";
        B <= "0011010110111010";
        C <= "0001110001000010";
        wait for clk_period;
        A <= "1111011010000101";
        B <= "1101100001110101";
        C <= "1110100011100000";
        wait for clk_period;
        A <= "0100000011101111";
        B <= "1111000010111110";
        C <= "1111010100001001";
        wait for clk_period;
        A <= "0000100100000111";
        B <= "0100100000001111";
        C <= "1000001100010101";
        wait for clk_period;
        A <= "1110110010100111";
        B <= "0010010110111101";
        C <= "0011000110100000";
        wait for clk_period;
        A <= "0111101101100010";
        B <= "1000100000101000";
        C <= "0110000111011000";
        wait for clk_period;
        A <= "1010010001101101";
        B <= "1101111101100110";
        C <= "0100100001010111";
        wait for clk_period;
        A <= "0100100011000111";
        B <= "1010110111111100";
        C <= "1110010110001011";
        wait for clk_period;
        A <= "1000000110101111";
        B <= "1100100001010010";
        C <= "1101111110010101";
        wait for clk_period;
        A <= "1110110001101111";
        B <= "1001100010011110";
        C <= "0101011001011111";
        wait for clk_period;
        A <= "1000110100001111";
        B <= "0110001100010100";
        C <= "0011111011000011";
        wait for clk_period;
        A <= "1101011100011110";
        B <= "0000010110011011";
        C <= "1011011100100110";
        wait for clk_period;
        A <= "0101011111100010";
        B <= "0010110101001011";
        C <= "1011011101010011";
        wait for clk_period;
        A <= "1100111111111111";
        B <= "0001111010001100";
        C <= "1100100011001101";
        wait for clk_period;
        A <= "1100100111000111";
        B <= "1111000111101001";
        C <= "1011001010011100";
        wait for clk_period;
        A <= "0010100110001100";
        B <= "0110111101000111";
        C <= "1010011001101100";
        wait for clk_period;
        A <= "0011010000010000";
        B <= "0011100111001101";
        C <= "0011001010101000";
        wait for clk_period;
        A <= "0101111000001000";
        B <= "0100110111100110";
        C <= "1011000111101111";
        wait for clk_period;
        A <= "1111110101111111";
        B <= "0001101101110000";
        C <= "0000001100110111";
        wait for clk_period;
        A <= "0100001101111111";
        B <= "1010100010110011";
        C <= "0100010100010100";
        wait for clk_period;
        A <= "1100000100001011";
        B <= "1000011100100110";
        C <= "0111010110101000";
        wait for clk_period;
        A <= "0000100010111111";
        B <= "1111111001010110";
        C <= "1110011010011010";
        wait for clk_period;
        A <= "1010111000000001";
        B <= "1001101100011001";
        C <= "0111111000010111";
        wait for clk_period;
        A <= "1011110000100000";
        B <= "0100011001110111";
        C <= "1000011001010000";
        wait for clk_period;
        A <= "1111000101000110";
        B <= "0100011010101100";
        C <= "0010110101100001";
        wait for clk_period;
        A <= "0010100100000100";
        B <= "1101100111011110";
        C <= "1011111000001010";
        wait for clk_period;
        A <= "1001010101001111";
        B <= "1101001101011111";
        C <= "1111110100111110";
        wait for clk_period;
        A <= "0101110111010110";
        B <= "1100011001000000";
        C <= "1110110111011101";
        wait for clk_period;
        A <= "0111011000101010";
        B <= "0001000101110111";
        C <= "0011111100010010";
        wait for clk_period;
        A <= "0100100100001011";
        B <= "1010001001110110";
        C <= "0011111101110011";
        wait for clk_period;
        A <= "0001101111011101";
        B <= "1101001110100110";
        C <= "1010100111101010";
        wait for clk_period;
        A <= "1110101101001001";
        B <= "1010000100001011";
        C <= "0001100010111010";
        wait for clk_period;
        A <= "1101101100100100";
        B <= "1010010000100000";
        C <= "0011001101001000";
        wait for clk_period;
        A <= "0110100111011111";
        B <= "0101100001000010";
        C <= "0001111010001110";
        wait for clk_period;
        A <= "1100111100111001";
        B <= "0010111111100000";
        C <= "0000110010010010";
        wait for clk_period;
        A <= "0000011011011000";
        B <= "1111111011011001";
        C <= "0011001111111000";
        wait for clk_period;
        A <= "0100100111100111";
        B <= "1101011001100001";
        C <= "1111000110111001";
        wait for clk_period;
        A <= "1100110000101111";
        B <= "1001010000011100";
        C <= "0001101100001011";
        wait for clk_period;
        A <= "0011010010111100";
        B <= "1100001111110010";
        C <= "0001001101000101";
        wait for clk_period;
        A <= "0101110100011101";
        B <= "0010110011101111";
        C <= "0000000011010110";
        wait for clk_period;
        A <= "1111011011111110";
        B <= "0110101100011110";
        C <= "0111011110000000";
        wait for clk_period;
        A <= "0100011000001110";
        B <= "1011110000000111";
        C <= "0101110001101100";
        wait for clk_period;
        A <= "1110101000011001";
        B <= "0010111001000100";
        C <= "0001100001011000";
        wait for clk_period;
        A <= "0010111100001011";
        B <= "1010011111100000";
        C <= "1111110010101111";
        wait for clk_period;
        A <= "0101000000001100";
        B <= "0000110010101000";
        C <= "1001010110011011";
        wait for clk_period;
        A <= "0101011110001010";
        B <= "1000010001010101";
        C <= "1111101001011111";
        wait for clk_period;
        A <= "0100000010010001";
        B <= "0101000011101011";
        C <= "0010001110111100";
        wait for clk_period;
        A <= "0010110011100110";
        B <= "1011111101000111";
        C <= "1101110001101101";
        wait for clk_period;
        A <= "1100110101101001";
        B <= "1100011010010100";
        C <= "1001101110110100";
        wait for clk_period;
        A <= "0000100000000000";
        B <= "1111001110111101";
        C <= "0011011100101111";
        wait for clk_period;
        A <= "1010110010000111";
        B <= "0010111011110001";
        C <= "0101101100100011";
        wait for clk_period;
        A <= "0000100010011010";
        B <= "1000100010010000";
        C <= "1111100000011010";
        wait for clk_period;
        A <= "1011010001110100";
        B <= "0101100010011011";
        C <= "1111010001000110";
        wait for clk_period;
        A <= "0101100001100010";
        B <= "1101111100110011";
        C <= "1011111001010000";
        wait for clk_period;
        A <= "1100011010110110";
        B <= "1001100101001010";
        C <= "0000000111011110";
        wait for clk_period;
        A <= "1110011101000111";
        B <= "0111100011111000";
        C <= "0010000110100111";
        wait for clk_period;
        A <= "0010101001011110";
        B <= "0011101011000011";
        C <= "0100110000001101";
        wait for clk_period;
        A <= "0001001100111111";
        B <= "0111111101111001";
        C <= "0010000110001000";
        wait for clk_period;
        A <= "0100110111000111";
        B <= "1011101101010101";
        C <= "1110001010010100";
        wait for clk_period;
        A <= "1000011011001001";
        B <= "1000011010010111";
        C <= "1001011011111010";
        wait for clk_period;
        A <= "0001111010101000";
        B <= "0010001000011011";
        C <= "1001011100000111";
        wait for clk_period;
        A <= "0001011001101101";
        B <= "1001100010011101";
        C <= "0011101101110000";
        wait for clk_period;
        A <= "1111001001000100";
        B <= "0010100100001011";
        C <= "1111111111010100";
        wait for clk_period;
        A <= "0100001000010111";
        B <= "1100011100101111";
        C <= "0000010010010111";
        wait for clk_period;
        A <= "1101101000100100";
        B <= "0001001100100010";
        C <= "0100100100000011";
        wait for clk_period;
        A <= "1000111100010010";
        B <= "0101110011100000";
        C <= "0010110010100110";
        wait for clk_period;
        A <= "0001111110100011";
        B <= "1001100100001001";
        C <= "1100011110100010";
        wait for clk_period;
        A <= "1101011000010101";
        B <= "1111111001111000";
        C <= "0111001000011111";
        wait for clk_period;
        A <= "1111001011101111";
        B <= "0000000011111110";
        C <= "0111111111010011";
        wait for clk_period;
        A <= "0000101001011111";
        B <= "0000111001101100";
        C <= "1010100100011100";
        wait for clk_period;
        A <= "1110101110111001";
        B <= "0101000101001110";
        C <= "1010101001000101";
        wait for clk_period;
        A <= "0000000111101101";
        B <= "0000000001111011";
        C <= "0100000000011001";
        wait for clk_period;
        A <= "0011100000000001";
        B <= "1100001100001001";
        C <= "0011011000000110";
        wait for clk_period;
        A <= "0000110010011110";
        B <= "1111100101010011";
        C <= "0111011010011011";
        wait for clk_period;
        A <= "1001011100010001";
        B <= "1011010111011000";
        C <= "0010000100110011";
        wait for clk_period;
        A <= "1011001001100111";
        B <= "1010011001001000";
        C <= "1100001110101011";
        wait for clk_period;
        A <= "1000100111110010";
        B <= "0101000111100110";
        C <= "0000100000100100";
        wait for clk_period;
        A <= "1011110110110011";
        B <= "1001101001100011";
        C <= "1100111101010101";
        wait for clk_period;
        A <= "0100100011000101";
        B <= "1001011100000010";
        C <= "1111001111111011";
        wait for clk_period;
        A <= "1001111111010000";
        B <= "1100001000110101";
        C <= "1100111000110010";
        wait for clk_period;
        A <= "1010111110000100";
        B <= "1111110101110101";
        C <= "1100110000010101";
        wait for clk_period;
        A <= "0111101011100101";
        B <= "1001100111111111";
        C <= "0101100010010111";
        wait for clk_period;
        A <= "1001110001111011";
        B <= "0011010011110000";
        C <= "1011110100011010";
        wait for clk_period;
        A <= "0100000110001100";
        B <= "0011011010110100";
        C <= "1101001111001110";
        wait for clk_period;
        A <= "1100101011100001";
        B <= "0011000110011001";
        C <= "1111010010010001";
        wait for clk_period;
        A <= "1000110101100111";
        B <= "1101100010111100";
        C <= "1101000001011001";
        wait for clk_period;
        A <= "1010001111111011";
        B <= "0100111100010101";
        C <= "1010001111000000";
        wait for clk_period;
        A <= "1011011111111111";
        B <= "0000110100110101";
        C <= "0010001011011001";
        wait for clk_period;
        A <= "0010010101001010";
        B <= "1010011011011100";
        C <= "0010110111111000";
        wait for clk_period;
        A <= "1111110111000110";
        B <= "1100000000010010";
        C <= "0100010011001110";
        wait for clk_period;
        A <= "0010001100001110";
        B <= "1011100011101000";
        C <= "1010110110110110";
        wait for clk_period;
        A <= "1010011000110110";
        B <= "0011100010011011";
        C <= "1000100000011011";
        wait for clk_period;
        A <= "1110110000000011";
        B <= "1110100100011010";
        C <= "1000011000100000";
        wait for clk_period;
        A <= "1110011010000011";
        B <= "1000000101000110";
        C <= "1110101000000001";
        wait for clk_period;
        A <= "0011010010100111";
        B <= "1000101110001111";
        C <= "1111010110100101";
        wait for clk_period;
        A <= "1011111001010110";
        B <= "1000111001111010";
        C <= "0010011010010001";
        wait for clk_period;
        A <= "0011010001011000";
        B <= "0110101100100001";
        C <= "1010001001001000";
        wait for clk_period;
        A <= "1001110111001000";
        B <= "1010100000010000";
        C <= "0000001100010101";
        wait for clk_period;
        A <= "1110011101001010";
        B <= "1111000000000011";
        C <= "0001010011110111";
        wait for clk_period;
        A <= "1100111110010100";
        B <= "1110100001011100";
        C <= "0110001110111111";
        wait for clk_period;
        A <= "1001010010010101";
        B <= "1111010010010001";
        C <= "1000110001100101";
        wait for clk_period;
        A <= "0000011010101000";
        B <= "0100100011110001";
        C <= "0011001000010111";
        wait for clk_period;
        A <= "1111001100111101";
        B <= "0001101101101100";
        C <= "1011111110111101";
        wait for clk_period;
        A <= "1100111001000100";
        B <= "0000000001011001";
        C <= "1011000010000001";
        wait for clk_period;
        A <= "0010110101001111";
        B <= "1010100010110101";
        C <= "0101110000111001";
        wait for clk_period;
        A <= "1011100100010011";
        B <= "1000100001101000";
        C <= "1101101001010110";
        wait for clk_period;
        A <= "0010110100000001";
        B <= "0100110001100011";
        C <= "1101111001010101";
        wait for clk_period;
        A <= "0000110100001111";
        B <= "0110110010010001";
        C <= "1001010110111101";
        wait for clk_period;
        A <= "0110110101111011";
        B <= "1101010110100100";
        C <= "0001111101110100";
        wait for clk_period;
        A <= "0000100101101011";
        B <= "0100111101101000";
        C <= "0000111110100010";
        wait for clk_period;
        A <= "0111110110100111";
        B <= "1001000110011010";
        C <= "1010111001001110";
        wait for clk_period;
        A <= "1111011000100111";
        B <= "1001101111011010";
        C <= "0011010110110101";
        wait for clk_period;
        A <= "0101100101110011";
        B <= "0100000011001100";
        C <= "1011010100110010";
        wait for clk_period;
        A <= "1011000111111010";
        B <= "1101010110111000";
        C <= "0010101000010000";
        wait for clk_period;
        A <= "1010001010000001";
        B <= "0100101001001110";
        C <= "1111011100110101";
        wait for clk_period;
        A <= "1001000001110010";
        B <= "0011101100110001";
        C <= "1101100111001001";
        wait for clk_period;
        A <= "0011101111100111";
        B <= "1010011111011100";
        C <= "1110011001100010";
        wait for clk_period;
        A <= "0101101000001100";
        B <= "1100110100101100";
        C <= "0110011001011000";
        wait for clk_period;
        A <= "0101111001101011";
        B <= "1111001110010000";
        C <= "1010111111001011";
        wait for clk_period;
        A <= "1101000000110101";
        B <= "0011010111001101";
        C <= "0111001111111100";
        wait for clk_period;
        A <= "0101100000101111";
        B <= "0010001111001111";
        C <= "0100011111001011";
        wait for clk_period;
        A <= "1001010001111011";
        B <= "0000111011000010";
        C <= "1000010100001001";
        wait for clk_period;
        A <= "1110000110011011";
        B <= "0100011010011100";
        C <= "0010011101101001";
        wait for clk_period;
        A <= "1101101110101010";
        B <= "1100100010100110";
        C <= "0110111110010001";
        wait for clk_period;
        A <= "0111010011100010";
        B <= "1001111101000000";
        C <= "1101100011100100";
        wait for clk_period;
        A <= "0110001000011000";
        B <= "1110110110100011";
        C <= "0000000000101011";
        wait for clk_period;
        A <= "0001100111111110";
        B <= "0011110111010011";
        C <= "1111111011110010";
        wait for clk_period;
        A <= "0010011011111000";
        B <= "1001000101100010";
        C <= "1101111100100011";
        wait for clk_period;
        A <= "1100100001001000";
        B <= "0111100001001000";
        C <= "1100100111000110";
        wait for clk_period;
        A <= "0100110101111000";
        B <= "1010001001111110";
        C <= "0011000010110010";
        wait for clk_period;
        A <= "1010000011011101";
        B <= "1111001011001100";
        C <= "1000110010110110";
        wait for clk_period;
        A <= "0110111100111001";
        B <= "0100010111001100";
        C <= "0010000101101110";
        wait for clk_period;
        A <= "1100011111110110";
        B <= "0100001100111110";
        C <= "1000001100110100";
        wait for clk_period;
        A <= "1101000000100001";
        B <= "1111100010001010";
        C <= "1010011001110001";
        wait for clk_period;
        A <= "1111110001000100";
        B <= "0110001000111011";
        C <= "1111100010011001";
        wait for clk_period;
        A <= "0001011100010001";
        B <= "1111101000101100";
        C <= "0011011001011100";
        wait for clk_period;
        A <= "0001111010001100";
        B <= "0110000111010001";
        C <= "1110100001101110";
        wait for clk_period;
        A <= "0000010000000111";
        B <= "1101111110111110";
        C <= "1010101001011000";
        wait for clk_period;
        A <= "1010101100001110";
        B <= "0001101000001101";
        C <= "1001110101001010";
        wait for clk_period;
        A <= "0100001110011111";
        B <= "1100000001110000";
        C <= "1011010111100010";
        wait for clk_period;
        A <= "1100001110111010";
        B <= "1010111100110000";
        C <= "0100001010000111";
        wait for clk_period;
        A <= "0000011000101101";
        B <= "1100101101001110";
        C <= "0111010111000100";
        wait for clk_period;
        A <= "0010110111110010";
        B <= "0000011111111011";
        C <= "0100010011110001";
        wait for clk_period;
        A <= "0101110001110001";
        B <= "0011110110101100";
        C <= "0010000100011011";
        wait for clk_period;
        A <= "0001111110110101";
        B <= "1011110010001000";
        C <= "0001001000010000";
        wait for clk_period;
        A <= "0110100100010110";
        B <= "0010001000110111";
        C <= "1100000100110111";
        wait for clk_period;
        A <= "0100011001011111";
        B <= "1001110000101000";
        C <= "0001000111000000";
        wait for clk_period;
        A <= "1100000000101001";
        B <= "0000011001101110";
        C <= "1000010011101000";
        wait for clk_period;
        A <= "0101111110110100";
        B <= "1001101001001011";
        C <= "0011000101010110";
        wait for clk_period;
        A <= "0010001001011100";
        B <= "1101110010000010";
        C <= "1010000001001100";
        wait for clk_period;
        A <= "0001101101101101";
        B <= "0100010110010101";
        C <= "0001010110001110";
        wait for clk_period;
        A <= "1001010011000001";
        B <= "0101111100010101";
        C <= "0001110100001011";
        wait for clk_period;
        A <= "1011110101101100";
        B <= "1100000111100101";
        C <= "1011111100000100";
        wait for clk_period;
        A <= "0111001101011001";
        B <= "1101111000100111";
        C <= "1010100110000011";
        wait for clk_period;
        A <= "0111110010101110";
        B <= "0100000011111010";
        C <= "0111010010011110";
        wait for clk_period;
        A <= "1001110111011100";
        B <= "0001011001110110";
        C <= "1010011101010100";
        wait for clk_period;
        A <= "1101011100011111";
        B <= "1101001101000011";
        C <= "0010001100000110";
        wait for clk_period;
        A <= "0010000100000111";
        B <= "1011111110111101";
        C <= "1101011111000111";
        wait for clk_period;
        A <= "1001100101000110";
        B <= "1100101001111001";
        C <= "1000010101011111";
        wait for clk_period;
        A <= "1111001011010100";
        B <= "0010010000010101";
        C <= "0101000111100100";
        wait for clk_period;
        A <= "0101011111011110";
        B <= "0000001111101001";
        C <= "0001100011101110";
        wait for clk_period;
        A <= "0100111000101000";
        B <= "0111111100011001";
        C <= "0010000100110011";
        wait for clk_period;
        A <= "0101000001000011";
        B <= "0110101100100100";
        C <= "0111111110100011";
        wait for clk_period;
        A <= "0010101101100010";
        B <= "0101010010011000";
        C <= "0000110111001001";
        wait for clk_period;
        A <= "0111111010110010";
        B <= "0011001111011101";
        C <= "0101010011000110";
        wait for clk_period;
        A <= "1000111011000001";
        B <= "1000100111100011";
        C <= "1010100111100100";
        wait for clk_period;
        A <= "0110101000100111";
        B <= "0000011010100000";
        C <= "1100011100111001";
        wait for clk_period;
        A <= "0011011000011110";
        B <= "0010010011110010";
        C <= "1011010101111111";
        wait for clk_period;
        A <= "1000000110110100";
        B <= "1111100001100110";
        C <= "0111110100101010";
        wait for clk_period;
        A <= "1010110000000010";
        B <= "0101101100010110";
        C <= "0010000100111001";
        wait for clk_period;
        A <= "1101010000011101";
        B <= "0000010101110111";
        C <= "0010110011010000";
        wait for clk_period;
        A <= "0111010010001101";
        B <= "0111001001000011";
        C <= "1001110110010011";
        wait for clk_period;
        A <= "1110010000000010";
        B <= "0110101011101111";
        C <= "0100111111001001";
        wait for clk_period;
        A <= "0101011111100010";
        B <= "0000101110100010";
        C <= "0001001001110101";
        wait for clk_period;
        A <= "1101001110100101";
        B <= "1011000101000011";
        C <= "0101001000011110";
        wait for clk_period;
        A <= "1001011010001110";
        B <= "1000100101011010";
        C <= "0111111110010010";
        wait for clk_period;
        A <= "0000110100101100";
        B <= "1001101101100110";
        C <= "0001110111111101";
        wait for clk_period;
        A <= "1011010111001000";
        B <= "0000001001000101";
        C <= "1111100100001010";
        wait for clk_period;
        A <= "0001011010110110";
        B <= "0110101101001001";
        C <= "1110110000000000";
        wait for clk_period;
        A <= "1101101101000001";
        B <= "1111000000001010";
        C <= "0101000000101111";
        wait for clk_period;
        A <= "1001010110011001";
        B <= "1100100011010101";
        C <= "1001000101001011";
        wait for clk_period;
        A <= "0001011101001100";
        B <= "0111001100110010";
        C <= "0010011010101001";
        wait for clk_period;
        A <= "1100000100010111";
        B <= "1010000001000101";
        C <= "1011000011111001";
        wait for clk_period;
        A <= "0101000100010111";
        B <= "0101010100100101";
        C <= "1110010101011011";
        wait for clk_period;
        A <= "0110000100111010";
        B <= "0110111110010010";
        C <= "0011100101100101";
        wait for clk_period;
        A <= "0001111010011111";
        B <= "0111110011001011";
        C <= "0101111000110010";
        wait for clk_period;
        A <= "1011010010011111";
        B <= "0011001111010110";
        C <= "0101101001101011";
        wait for clk_period;
        A <= "1111010010001110";
        B <= "1000100101111011";
        C <= "1100001101011011";
        wait for clk_period;
        A <= "1010001100010111";
        B <= "0101110000000010";
        C <= "0001111010110100";
        wait for clk_period;
        A <= "1111011010100010";
        B <= "1100110100000101";
        C <= "1111010011101101";
        wait for clk_period;
        A <= "1111110111010000";
        B <= "1010001100010010";
        C <= "0001011000101011";
        wait for clk_period;
        A <= "0111111001001100";
        B <= "1000101011111111";
        C <= "1001100000111000";
        wait for clk_period;
        A <= "1001111100110011";
        B <= "1100011111011001";
        C <= "1100010100011101";
        wait for clk_period;
        A <= "0001000100111111";
        B <= "0000000111111101";
        C <= "0011100100111001";
        wait for clk_period;
        A <= "1101011111001000";
        B <= "1101011001101100";
        C <= "0110010110110110";
        wait for clk_period;
        A <= "1000010000100001";
        B <= "0101111111011010";
        C <= "0111011011011011";
        wait for clk_period;
        A <= "1011111110000011";
        B <= "0101100110101000";
        C <= "0100010111111111";
        wait for clk_period;
        A <= "1101010001011001";
        B <= "0010111001010001";
        C <= "1110100110101001";
        wait for clk_period;
        A <= "1011000101100111";
        B <= "0110000000110000";
        C <= "1111010001000000";
        wait for clk_period;
        A <= "1100000111011101";
        B <= "0110000100011000";
        C <= "1100111111100010";
        wait for clk_period;
        A <= "1110000011000111";
        B <= "0110100011111111";
        C <= "1100000000101101";
        wait for clk_period;
        A <= "0000010011101110";
        B <= "1101101011111110";
        C <= "1011011011001010";
        wait for clk_period;
        A <= "1011110000110000";
        B <= "0011001011001110";
        C <= "1111011110000110";
        wait for clk_period;
        A <= "1110010001110000";
        B <= "1100001001010011";
        C <= "1001011000101110";
        wait for clk_period;
        A <= "1101000111111100";
        B <= "1101011011111110";
        C <= "0110101110101101";
        wait for clk_period;
        A <= "0100011100011100";
        B <= "0111011110101110";
        C <= "1010100110011011";
        wait for clk_period;
        A <= "1101010001010111";
        B <= "0101101011000000";
        C <= "0000010000000000";
        wait for clk_period;
        A <= "1000011011101011";
        B <= "1110111001000100";
        C <= "1000101010101011";
        wait for clk_period;
        A <= "0000010000001111";
        B <= "1100111110101001";
        C <= "1110110101000011";
        wait for clk_period;
        A <= "0101100001010100";
        B <= "0110010111100010";
        C <= "1000001010000001";
        wait for clk_period;
        A <= "0010101110100001";
        B <= "1111101100001010";
        C <= "0100010101100001";
        wait for clk_period;
        A <= "1101010001110000";
        B <= "1111100101110001";
        C <= "1001000110101010";
        wait for clk_period;
        A <= "1100101110101011";
        B <= "0000000101101000";
        C <= "0111010010111001";
        wait for clk_period;
        A <= "0101000110101111";
        B <= "1111110100010111";
        C <= "0110100100100010";
        wait for clk_period;
        A <= "0000101010011100";
        B <= "1001101010100100";
        C <= "0100010101110011";
        wait for clk_period;
        A <= "0100011000101001";
        B <= "0011001100011000";
        C <= "1001000001011001";
        wait for clk_period;
        A <= "0101010110101111";
        B <= "1010010001111100";
        C <= "1001100100100001";
        wait for clk_period;
        A <= "1011111101010010";
        B <= "1111111001001011";
        C <= "1100001010101111";
        wait for clk_period;
        A <= "1001100111010011";
        B <= "1011011110011111";
        C <= "0101100100000001";
        wait for clk_period;
        A <= "1000111101010100";
        B <= "1010000011010110";
        C <= "1011000000000010";
        wait for clk_period;
        A <= "1111111110011101";
        B <= "0011010100111000";
        C <= "0000010100110010";
        wait for clk_period;
        A <= "1010010000001110";
        B <= "0101101000001111";
        C <= "0011111010110111";
        wait for clk_period;
        A <= "1001111000101110";
        B <= "1010111100000000";
        C <= "0110111110001010";
        wait for clk_period;
        A <= "0010111011110001";
        B <= "0101000111001000";
        C <= "0110100100100010";
        wait for clk_period;
        A <= "0001011100100100";
        B <= "1001101000001110";
        C <= "1111100000110011";
        wait for clk_period;
        A <= "0110010110111010";
        B <= "0110101010110110";
        C <= "0011000000110000";
        wait for clk_period;
        A <= "0011000010001001";
        B <= "0011111110001011";
        C <= "0000001000010011";
        wait for clk_period;
        A <= "1001101110001010";
        B <= "0111000110010100";
        C <= "0100011000010001";
        wait for clk_period;
        A <= "1000010000111001";
        B <= "0111000111000011";
        C <= "1000111100100101";
        wait for clk_period;
        A <= "1111011010001110";
        B <= "0101100011001011";
        C <= "1110101001101000";
        wait for clk_period;
        A <= "1110110001100101";
        B <= "0001101110110100";
        C <= "0110111111001000";
        wait for clk_period;
        A <= "0111001110010011";
        B <= "1000101011100100";
        C <= "0101001111101100";
        wait for clk_period;
        A <= "1110000100101001";
        B <= "0111100011111000";
        C <= "0011101101001000";
        wait for clk_period;
        A <= "1110010100111010";
        B <= "0000011111101011";
        C <= "1010001000001011";
        wait for clk_period;
        A <= "1011000011100000";
        B <= "0011110001100110";
        C <= "0110001110000010";
        wait for clk_period;
        A <= "1101111000101110";
        B <= "0110000010001111";
        C <= "0111010011101010";
        wait for clk_period;
        A <= "0100010101100011";
        B <= "1110111010001101";
        C <= "1000000001011100";
        wait for clk_period;
        A <= "0101000010101000";
        B <= "1001001011110100";
        C <= "0101100000001111";
        wait for clk_period;
        A <= "1000101110000110";
        B <= "0110000000001110";
        C <= "1111100000111010";
        wait for clk_period;
        A <= "1001100110100110";
        B <= "1101111110101111";
        C <= "1111100011100010";
        wait for clk_period;
        A <= "0101101101000000";
        B <= "1111000111100110";
        C <= "0001111000110011";
        wait for clk_period;
        A <= "0101001100001101";
        B <= "0110110101010011";
        C <= "1010011111010101";
        wait for clk_period;
        A <= "1011100010011111";
        B <= "1000111011110000";
        C <= "1000111111101111";
        wait for clk_period;
        A <= "0101011011101101";
        B <= "0011101001100011";
        C <= "1110101001000100";
        wait for clk_period;
        A <= "1010001010000010";
        B <= "1110110000000001";
        C <= "0110110000110011";
        wait for clk_period;
        A <= "1010101010001010";
        B <= "1010111101001111";
        C <= "0111010001101010";
        wait for clk_period;
        A <= "0011110100011100";
        B <= "1011100101000011";
        C <= "0001001101110101";
        wait for clk_period;
        A <= "0001010100100011";
        B <= "0010010000110100";
        C <= "1010100101111000";
        wait for clk_period;
        A <= "1001100000000010";
        B <= "1110010010111101";
        C <= "1010110010111101";
        wait for clk_period;
        A <= "0110000000011111";
        B <= "0101110001100100";
        C <= "0101110011010110";
        wait for clk_period;
        A <= "0111010000110100";
        B <= "0101011110010000";
        C <= "0110001010001010";
        wait for clk_period;
        A <= "1100010111101001";
        B <= "1001000101100101";
        C <= "1001011101011111";
        wait for clk_period;
        A <= "1010011001000101";
        B <= "0000010110001000";
        C <= "1110000101110001";
        wait for clk_period;
        A <= "1000001001010010";
        B <= "1100100111000010";
        C <= "1010111110001111";
        wait for clk_period;
        A <= "0111111010100100";
        B <= "0000011010011111";
        C <= "1101010011010111";
        wait for clk_period;
        A <= "0011100101001101";
        B <= "0100011101000001";
        C <= "1110000011100100";
        wait for clk_period;
        A <= "0110101101100011";
        B <= "0011001000100100";
        C <= "1100110011100001";
        wait for clk_period;
        A <= "0100101110011000";
        B <= "1110111101011110";
        C <= "1100001000011100";
        wait for clk_period;
        A <= "0000100110111000";
        B <= "1010101000010111";
        C <= "0101001100111110";
        wait for clk_period;
        A <= "1100111111101001";
        B <= "0011011001001100";
        C <= "1000110101101010";
        wait for clk_period;
        A <= "0000000100011000";
        B <= "1110100111111111";
        C <= "1111010001000010";
        wait for clk_period;
        A <= "0010010110000110";
        B <= "1110010111101000";
        C <= "0111011110101111";
        wait for clk_period;
        A <= "0100010111110010";
        B <= "1010110001111001";
        C <= "1010110100101111";
        wait for clk_period;
        A <= "1101011101001000";
        B <= "0001011111001100";
        C <= "0111001101100101";
        wait for clk_period;
        A <= "1100001011010101";
        B <= "1001111011000000";
        C <= "1101000101000100";
        wait for clk_period;
        A <= "1110111000111110";
        B <= "0110111111110010";
        C <= "1101011011000001";
        wait for clk_period;
        A <= "1001111011001111";
        B <= "0110101101001010";
        C <= "1010110111110010";
        wait for clk_period;
        A <= "1000110011010000";
        B <= "0010111001011010";
        C <= "0011110100110110";
        wait for clk_period;
        A <= "1110110110111000";
        B <= "0010010101001101";
        C <= "1100100011111110";
        wait for clk_period;
        A <= "0110100010010110";
        B <= "1101110111100011";
        C <= "0110110110010000";
        wait for clk_period;
        A <= "1100000011110100";
        B <= "1001110111100000";
        C <= "0010011000010110";
        wait for clk_period;
        A <= "0011111010001011";
        B <= "0111011000001010";
        C <= "1110111011110010";
        wait for clk_period;
        A <= "1000100011111111";
        B <= "1100100111100100";
        C <= "1010111101101000";
        wait for clk_period;
        A <= "0101000100011001";
        B <= "1100110001101101";
        C <= "1100010111001111";
        wait for clk_period;
        A <= "0100110110111100";
        B <= "1100001110100000";
        C <= "1011100101001011";
        wait for clk_period;
        A <= "0111011110111110";
        B <= "0000000011100110";
        C <= "1101100100000011";
        wait for clk_period;
        A <= "0110101101100001";
        B <= "1110011010011000";
        C <= "0101000011001101";
        wait for clk_period;
        A <= "1000110011101011";
        B <= "1010100101001110";
        C <= "1010000111100010";
        wait for clk_period;
        A <= "1101010010111010";
        B <= "1100001010010011";
        C <= "0000011111110111";
        wait for clk_period;
        A <= "1011000011001110";
        B <= "1001000111100011";
        C <= "1001000100101111";
        wait for clk_period;
        A <= "0010101010110000";
        B <= "0001110001000111";
        C <= "1111011000010100";
        wait for clk_period;
        A <= "0101111110011110";
        B <= "0100101100111011";
        C <= "0001111000001111";
        wait for clk_period;
        A <= "0101010111011001";
        B <= "0010001110000011";
        C <= "0100110101010101";
        wait for clk_period;
        A <= "0011101110010101";
        B <= "1000111110000000";
        C <= "1101010011101101";
        wait for clk_period;
        A <= "1101001100111000";
        B <= "0000111010011011";
        C <= "1101101000111100";
        wait for clk_period;
        A <= "1000110101100100";
        B <= "0010001010100110";
        C <= "1001010110110010";
        wait for clk_period;
        A <= "0010111111000010";
        B <= "1110101000110110";
        C <= "1001010010111110";
        wait for clk_period;
        A <= "0000111000110000";
        B <= "0110111101001111";
        C <= "0011001101000100";
        wait for clk_period;
        A <= "0010110001011111";
        B <= "0111010101100101";
        C <= "0001110111011100";
        wait for clk_period;
        A <= "0011000000000101";
        B <= "0110001011001011";
        C <= "1001110000001000";
        wait for clk_period;
        A <= "0111110101001000";
        B <= "0011111101010101";
        C <= "0000101000100011";
        wait for clk_period;
        A <= "0010011111110000";
        B <= "0111001101110100";
        C <= "1100010001010010";
        wait for clk_period;
        A <= "0011100011000100";
        B <= "0100111101101001";
        C <= "0111001010110011";
        wait for clk_period;
        A <= "1100110100111101";
        B <= "0101011101100101";
        C <= "0011101111101010";
        wait for clk_period;
        A <= "1010010101001100";
        B <= "0110010011000011";
        C <= "0010000101001010";
        wait for clk_period;
        A <= "0000011000011001";
        B <= "0001001000010111";
        C <= "1001100111011100";
        wait for clk_period;
        A <= "0100000101110001";
        B <= "1101111111110101";
        C <= "0010011000100111";
        wait for clk_period;
        A <= "0001000111001110";
        B <= "0111011110010110";
        C <= "1100001101111010";
        wait for clk_period;
        A <= "0110000001101011";
        B <= "1111101010000010";
        C <= "0000000111010101";
        wait for clk_period;
        A <= "0100101000100100";
        B <= "1100111010101010";
        C <= "1001101110100001";
        wait for clk_period;
        A <= "0011000000110100";
        B <= "1110111011101001";
        C <= "1000111011110110";
        wait for clk_period;
        A <= "1010011000010110";
        B <= "0110110110011110";
        C <= "1010011100011010";
        wait for clk_period;
        A <= "1000101001100001";
        B <= "1100111111100110";
        C <= "0001111001101111";
        wait for clk_period;
        A <= "1100000111101010";
        B <= "0111100100101010";
        C <= "0101011110011110";
        wait for clk_period;
        A <= "1001000001110010";
        B <= "1000001000111001";
        C <= "0100001001101100";
        wait for clk_period;
        A <= "0101011001000010";
        B <= "1111010000001100";
        C <= "1101000010111001";
        wait for clk_period;
        A <= "0001101110110001";
        B <= "0110111110110000";
        C <= "1110100100100100";
        wait for clk_period;
        A <= "0001000001101001";
        B <= "1101010010000000";
        C <= "1110100101011011";
        wait for clk_period;
        A <= "0000011100011100";
        B <= "1000100011010000";
        C <= "1011011001001111";
        wait for clk_period;
        A <= "0110100100010111";
        B <= "0010100001100101";
        C <= "1000110111011011";
        wait for clk_period;
        A <= "1101000010111000";
        B <= "0000100010000000";
        C <= "0000001011100011";
        wait for clk_period;
        A <= "0011010001110001";
        B <= "0001100111000001";
        C <= "1001100001011100";
        wait for clk_period;
        A <= "1110100110101111";
        B <= "0010001011000101";
        C <= "1011100010111101";
        wait for clk_period;
        A <= "1010000001100101";
        B <= "0000011110000101";
        C <= "0111010101001111";
        wait for clk_period;
        A <= "1100111110011101";
        B <= "1101101001101111";
        C <= "1010111111110001";
        wait for clk_period;
        A <= "0100110101010000";
        B <= "1110111010000001";
        C <= "0111111101001101";
        wait for clk_period;
        A <= "0010001101100000";
        B <= "1000010010101111";
        C <= "1110001100100111";
        wait for clk_period;
        A <= "0011101111101000";
        B <= "0010011101100111";
        C <= "1001011101011000";
        wait for clk_period;
        A <= "0000010101011010";
        B <= "1011111011110011";
        C <= "1110100000010001";
        wait for clk_period;
        A <= "1110001001011001";
        B <= "1110010000111001";
        C <= "0000110110011100";
        wait for clk_period;
        A <= "1000101000000010";
        B <= "0111011101011110";
        C <= "1000101000010010";
        wait for clk_period;
        A <= "0111001000100110";
        B <= "1010010001011000";
        C <= "1110001111001000";
        wait for clk_period;
        A <= "1110101101010010";
        B <= "1100111000100111";
        C <= "1110011110100001";
        wait for clk_period;
        A <= "0110111001110101";
        B <= "0001101000110010";
        C <= "0100110000000010";
        wait for clk_period;
        A <= "1101011000011011";
        B <= "0110010001001111";
        C <= "0011101001000011";
        wait for clk_period;
        A <= "1111001001110110";
        B <= "0110010111000011";
        C <= "1001101011001000";
        wait for clk_period;
        A <= "1001101100111010";
        B <= "1110101010111110";
        C <= "0111000000010011";
        wait for clk_period;
        A <= "1101000000101111";
        B <= "0110101110100110";
        C <= "0000010000110010";
        wait for clk_period;
        A <= "1101001011101101";
        B <= "0011110100110100";
        C <= "1101111100010110";
        wait for clk_period;
        A <= "0011011110010110";
        B <= "0000001100111110";
        C <= "1000000110011100";
        wait for clk_period;
        A <= "0000110101010010";
        B <= "0101011010111011";
        C <= "0111110000010101";
        wait for clk_period;
        A <= "0010011001110100";
        B <= "0000000111001111";
        C <= "1110100000010110";
        wait for clk_period;
        A <= "1000110000011101";
        B <= "0001100100111000";
        C <= "0011011111100000";
        wait for clk_period;
        A <= "1100101001011011";
        B <= "0111011100101001";
        C <= "0110000110110110";
        wait for clk_period;
        A <= "1100101110101010";
        B <= "1010000000101111";
        C <= "0111111011110000";
        wait for clk_period;
        A <= "0001010011101011";
        B <= "0111000000111000";
        C <= "1101000000011000";
        wait for clk_period;
        A <= "1110011010001001";
        B <= "0100010011010101";
        C <= "0001111001111110";
        wait for clk_period;
        A <= "1000010111111011";
        B <= "1011101100011000";
        C <= "1000101101000000";
        wait for clk_period;
        A <= "0010100001001001";
        B <= "1111101100100111";
        C <= "0100011111001111";
        wait for clk_period;
        A <= "0001010011110010";
        B <= "1010000001111001";
        C <= "1010100001110100";
        wait for clk_period;
        A <= "0011110000101000";
        B <= "0111101001110010";
        C <= "0111110010100001";
        wait for clk_period;
        A <= "1110100111111010";
        B <= "1011100011000010";
        C <= "1101000010100111";
        wait for clk_period;
        A <= "1000001101101000";
        B <= "0100000010110010";
        C <= "0001101111110001";
        wait for clk_period;
        A <= "0111100001100100";
        B <= "1001101100110000";
        C <= "0001110111001001";
        wait for clk_period;
        A <= "0001101010011010";
        B <= "1010000111100011";
        C <= "0100001110000111";
        wait for clk_period;
        A <= "1111011100100101";
        B <= "1011000010110111";
        C <= "0010100010100111";
        wait for clk_period;
        A <= "1001100001100000";
        B <= "1001101111110100";
        C <= "0101000100111000";
        wait for clk_period;
        A <= "0011110111000001";
        B <= "1111001110010011";
        C <= "0001010010100100";
        wait for clk_period;
        A <= "1001000101110101";
        B <= "0010101000111001";
        C <= "1101100000100110";
        wait for clk_period;
        A <= "0110110000110010";
        B <= "1110111101100101";
        C <= "1010011001011111";
        wait for clk_period;
        A <= "1001000110011000";
        B <= "1000111100011110";
        C <= "0111100001010101";
        wait for clk_period;
        A <= "0001001100111011";
        B <= "1001100011101110";
        C <= "0000110110000100";
        wait for clk_period;
        A <= "1001001011000010";
        B <= "1011010111101111";
        C <= "0010001001010101";
        wait for clk_period;
        A <= "0011100000010110";
        B <= "0001101110011111";
        C <= "1101011001001101";
        wait for clk_period;
        A <= "1111111111010100";
        B <= "1000001010010100";
        C <= "0001001101100000";
        wait for clk_period;
        A <= "1101001001011000";
        B <= "0001000101101011";
        C <= "1010100000010100";
        wait for clk_period;
        A <= "1000110100100011";
        B <= "0010111001001101";
        C <= "1101110001000110";
        wait for clk_period;
        A <= "0000110111001110";
        B <= "1111100000100011";
        C <= "0111011111010110";
        wait for clk_period;
        A <= "1111111110111011";
        B <= "1110100110111111";
        C <= "0001101010101101";
        wait for clk_period;
        A <= "1111010101011010";
        B <= "0110000011111001";
        C <= "0101001001000000";
        wait for clk_period;
        A <= "0001110010011101";
        B <= "1101011011111100";
        C <= "0111110000111100";
        wait for clk_period;
        A <= "0011010111101101";
        B <= "0110001011000000";
        C <= "1001110101001011";
        wait for clk_period;
        A <= "1011101000111010";
        B <= "1001000100001101";
        C <= "0101101101000100";
        wait for clk_period;
        A <= "0101010010110000";
        B <= "1001100110010110";
        C <= "1111101100000011";
        wait for clk_period;
        A <= "1000001101010000";
        B <= "0011010010010001";
        C <= "1110000111000100";
        wait for clk_period;
        A <= "1011000101000000";
        B <= "1011000110000111";
        C <= "1100000010010110";
        wait for clk_period;
        A <= "1001100111001010";
        B <= "1101010010001111";
        C <= "1010100100011000";
        wait for clk_period;
        A <= "1000111010110010";
        B <= "1011101100000000";
        C <= "0100010011010100";
        wait for clk_period;
        A <= "1100010100000011";
        B <= "1010001111111100";
        C <= "1110111001010110";
        wait for clk_period;
        A <= "0111010001010110";
        B <= "1000101011110100";
        C <= "0100110001011110";
        wait for clk_period;
        A <= "1001111111010110";
        B <= "0000100001110011";
        C <= "1000110101001100";
        wait for clk_period;
        A <= "0110100101000110";
        B <= "1110100000000111";
        C <= "0010110000110111";
        wait for clk_period;
        A <= "1011101111110100";
        B <= "0000001110011110";
        C <= "0110001101000101";
        wait for clk_period;
        A <= "1111110000101011";
        B <= "0110110111100011";
        C <= "1101011111101100";
        wait for clk_period;
        A <= "1000010100111110";
        B <= "1010010110000111";
        C <= "1100100100100110";
        wait for clk_period;
        A <= "1011011001010001";
        B <= "1010100100000100";
        C <= "1101100001101110";
        wait for clk_period;
        A <= "1010011011111100";
        B <= "0010110111001001";
        C <= "0001110000000011";
        wait for clk_period;
        A <= "0110011000011011";
        B <= "0110111101011011";
        C <= "0011110100101010";
        wait for clk_period;
        A <= "0010110001100010";
        B <= "1010110001011001";
        C <= "1010110111110100";
        wait for clk_period;
        A <= "1001110100100111";
        B <= "1110111100010001";
        C <= "1010100010011111";
        wait for clk_period;
        A <= "0011001101111010";
        B <= "0110100001001000";
        C <= "1101101111110101";
        wait for clk_period;
        A <= "0001010100110110";
        B <= "0011010011011100";
        C <= "1011111010100001";
        wait for clk_period;
        A <= "1011011001000011";
        B <= "1010011000100100";
        C <= "0011000011100001";
        wait for clk_period;
        A <= "0100001110001000";
        B <= "0111100000011001";
        C <= "0100011001101010";
        wait for clk_period;
        A <= "1111100110010101";
        B <= "0100100001000110";
        C <= "0000001110100011";
        wait for clk_period;
        A <= "1101010100001010";
        B <= "0100110111001001";
        C <= "0000110010001000";
        wait for clk_period;
        A <= "0010010100100011";
        B <= "0101001111011111";
        C <= "1010011110111011";
        wait for clk_period;
        A <= "0100110001011011";
        B <= "1000100011101011";
        C <= "0010100101011000";
        wait for clk_period;
        A <= "1001000110111110";
        B <= "0111001011100011";
        C <= "0100010110010101";
        wait for clk_period;
        A <= "1110111111001001";
        B <= "1100010110101010";
        C <= "0010101111011000";
        wait for clk_period;
        A <= "1100011111011100";
        B <= "0000111011000001";
        C <= "0100001111111100";
        wait for clk_period;
        A <= "1011101100011000";
        B <= "0101011011001010";
        C <= "0110110101010001";
        wait for clk_period;
        A <= "0001010011100110";
        B <= "1010001111101000";
        C <= "0001101110011110";
        wait for clk_period;
        A <= "0001000110101000";
        B <= "0101001011000110";
        C <= "0100011100000000";
        wait for clk_period;
        A <= "0011001000100101";
        B <= "1001011000001001";
        C <= "0100001001110110";
        wait for clk_period;
        A <= "1100101010011010";
        B <= "1101010111011101";
        C <= "1001001100111000";
        wait for clk_period;
        A <= "1110000001111001";
        B <= "0101000111001011";
        C <= "1101110100001010";
        wait for clk_period;
        A <= "1010000011110110";
        B <= "1001100000101101";
        C <= "0000011101001110";
        wait for clk_period;
        A <= "0011110010110011";
        B <= "0101110010001100";
        C <= "1110010110100011";
        wait for clk_period;
        A <= "0100100110110011";
        B <= "1101011010010100";
        C <= "0111101111111100";
        wait for clk_period;
        A <= "0010011011111101";
        B <= "0010111011101010";
        C <= "1011101110100001";
        wait for clk_period;
        A <= "1101010000000010";
        B <= "0101011010111101";
        C <= "0111011000111010";
        wait for clk_period;
        A <= "0011111001000001";
        B <= "0100100011001001";
        C <= "0000111100010100";
        wait for clk_period;
        A <= "1110000110001110";
        B <= "0111011010100011";
        C <= "0100010100011010";
        wait for clk_period;
        A <= "0111111010001010";
        B <= "0011100101001001";
        C <= "0010011010110000";
        wait for clk_period;
        A <= "0010000100100011";
        B <= "1011011111001000";
        C <= "0010010011100010";
        wait for clk_period;
        A <= "1010110011110100";
        B <= "0100110010100111";
        C <= "1101000101011010";
        wait for clk_period;
        A <= "1101010100000000";
        B <= "0100000000011001";
        C <= "0010101101010001";
        wait for clk_period;
        A <= "0010001100000010";
        B <= "0111011100000001";
        C <= "1110111100001000";
        wait for clk_period;
        A <= "0000101000000110";
        B <= "1001100000001110";
        C <= "0010100101110001";
        wait for clk_period;
        A <= "0100001101000110";
        B <= "0001010001010110";
        C <= "1001010110000010";
        wait for clk_period;
        A <= "0110010001100011";
        B <= "1000101001100011";
        C <= "1001110110001011";
        wait for clk_period;
        A <= "1100111000011010";
        B <= "1011000010011100";
        C <= "1110111010101011";
        wait for clk_period;
        A <= "0100000000111000";
        B <= "1100101010101101";
        C <= "1111100000010011";
        wait for clk_period;
        A <= "1001101111010111";
        B <= "0010010011001110";
        C <= "1101110000101110";
        wait for clk_period;
        A <= "1100100100101100";
        B <= "1001111010110101";
        C <= "1001001010011011";
        wait for clk_period;
        A <= "1101100111110011";
        B <= "0001111110100110";
        C <= "0111001101011011";
        wait for clk_period;
        A <= "0111011001001001";
        B <= "0110100010100010";
        C <= "0111100000101001";
        wait for clk_period;
        A <= "0010010011011111";
        B <= "0000000100100101";
        C <= "0010101010000001";
        wait for clk_period;
        A <= "1000000110101100";
        B <= "1011001110101101";
        C <= "1001111000011010";
        wait for clk_period;
        A <= "0101111101001110";
        B <= "1101010010101100";
        C <= "0010101000111101";
        wait for clk_period;
        A <= "0101110001000000";
        B <= "1111000110010101";
        C <= "0100000100011110";
        wait for clk_period;
        A <= "0111101011000001";
        B <= "1000000100111111";
        C <= "0000101010001001";
        wait for clk_period;
        A <= "0010010110011111";
        B <= "1111101010010100";
        C <= "1111111001111001";
        wait for clk_period;
        A <= "0110000011000010";
        B <= "0100011101011100";
        C <= "0111011010010000";
        wait for clk_period;
        A <= "0010010000000001";
        B <= "0101001000001011";
        C <= "1101110110100011";
        wait for clk_period;
        A <= "0011000111101010";
        B <= "1111001010110011";
        C <= "0011001100100101";
        wait for clk_period;
        A <= "0111110010100100";
        B <= "0001111010010011";
        C <= "0011000111111000";
        wait for clk_period;
        A <= "0110001001001000";
        B <= "0110011100111010";
        C <= "0011110011101101";
        wait for clk_period;
        A <= "1000101101100100";
        B <= "1000000110111000";
        C <= "0010110001101111";
        wait for clk_period;
        A <= "0100010001000011";
        B <= "0110111011011010";
        C <= "0100101010011011";
        wait for clk_period;
        A <= "0100010101011000";
        B <= "0010111111011111";
        C <= "1111011000101111";
        wait for clk_period;
        A <= "0111111001011101";
        B <= "1110001100110010";
        C <= "1010001111101011";
        wait for clk_period;
        A <= "0000010100110011";
        B <= "0001001000110011";
        C <= "0111110000001111";
        wait for clk_period;
        A <= "1001111010111111";
        B <= "0010001100100001";
        C <= "1110101010001110";
        wait for clk_period;
        A <= "1010100011100111";
        B <= "1000001001001111";
        C <= "1101100110100011";
        wait for clk_period;
        A <= "0010010110000111";
        B <= "0010011110101010";
        C <= "0001011000111010";
        wait for clk_period;
        A <= "1010110000111011";
        B <= "0000001110100101";
        C <= "0101010110011000";
        wait for clk_period;
        A <= "1011010011100001";
        B <= "1000110001100100";
        C <= "0101111010111001";
        wait for clk_period;
        A <= "1100010111010100";
        B <= "1010001110101011";
        C <= "0001001000001100";
        wait for clk_period;
        A <= "0011101000010100";
        B <= "0110110111011110";
        C <= "0011101011010101";
        wait for clk_period;
        A <= "0001001010111111";
        B <= "0011010101101011";
        C <= "1010101000100111";
        wait for clk_period;
        A <= "0111011011000110";
        B <= "0000100110110110";
        C <= "0001000111001011";
        wait for clk_period;
        A <= "1001111001010101";
        B <= "0111110110101100";
        C <= "0111010001001101";
        wait for clk_period;
        A <= "0001100000110001";
        B <= "0001000001101011";
        C <= "0100011001101100";
        wait for clk_period;
        A <= "1110101110010110";
        B <= "0110110001010010";
        C <= "1101110110000111";
        wait for clk_period;
        A <= "0111101111011101";
        B <= "1101001101100011";
        C <= "1101110100001111";
        wait for clk_period;
        A <= "1100100100110000";
        B <= "0000110110101011";
        C <= "0010000010111101";
        wait for clk_period;
        A <= "1000111100101001";
        B <= "0111010111110011";
        C <= "1011111010101111";
        wait for clk_period;
        A <= "1110110110010101";
        B <= "0011010010011001";
        C <= "1110101100011101";
        wait for clk_period;
        A <= "1000101001111001";
        B <= "1111101010110101";
        C <= "1010100101010111";
        wait for clk_period;
        A <= "1110010100000011";
        B <= "1000000000000110";
        C <= "0000010001100000";
        wait for clk_period;
        A <= "1101010010000011";
        B <= "0000101111011110";
        C <= "1000101100011101";
        wait for clk_period;
        A <= "0001010010111001";
        B <= "0100101011101100";
        C <= "0001000001010100";
        wait for clk_period;
        A <= "0101110111101110";
        B <= "0011101001000001";
        C <= "1001110001011010";
        wait for clk_period;
        A <= "1010000001011001";
        B <= "0100000010001000";
        C <= "0000010110001011";
        wait for clk_period;
        A <= "0000111011011001";
        B <= "0000001111010100";
        C <= "0100101001011110";
        wait for clk_period;
        A <= "1010001111001011";
        B <= "0101010011000110";
        C <= "1110011101001001";
        wait for clk_period;
        A <= "1100110111110000";
        B <= "1100010101010101";
        C <= "1100110000111110";
        wait for clk_period;
        A <= "1010111010010011";
        B <= "1100010111110110";
        C <= "0000101110011001";
        wait for clk_period;
        A <= "0011100000010100";
        B <= "1000000100110011";
        C <= "1011011001001110";
        wait for clk_period;
        A <= "1011110011001101";
        B <= "1111111001010111";
        C <= "0110110111001011";
        wait for clk_period;
        A <= "0111000101110111";
        B <= "0110101100011110";
        C <= "0011101100110001";
        wait for clk_period;
        A <= "1011010101101010";
        B <= "1000101010011101";
        C <= "1111011111100000";
        wait for clk_period;
        A <= "1101001111001111";
        B <= "1111100001110111";
        C <= "1111101101111110";
        wait for clk_period;
        A <= "0010001010111111";
        B <= "1101000100001111";
        C <= "0000011000011110";
        wait for clk_period;
        A <= "0101000010001000";
        B <= "0001000101100011";
        C <= "0100100111010101";
        wait for clk_period;
        A <= "1010101001010100";
        B <= "0111001011101111";
        C <= "1110011010100100";
        wait for clk_period;
        A <= "0100100011111001";
        B <= "0010001101101110";
        C <= "1101111001100100";
        wait for clk_period;
        A <= "1100111010001000";
        B <= "1001010000110010";
        C <= "0011110110100100";
        wait for clk_period;
        A <= "0011011110101011";
        B <= "1110001011011110";
        C <= "1100111111101011";
        wait for clk_period;
        A <= "0110111011100011";
        B <= "0010001110100100";
        C <= "1010010101110000";
        wait for clk_period;
        A <= "0100101111100100";
        B <= "1110011111110011";
        C <= "0111001001101010";
        wait for clk_period;
        A <= "0001000010000011";
        B <= "0110001110011010";
        C <= "1001011111110011";
        wait for clk_period;
        A <= "1111011100001000";
        B <= "0011011010001111";
        C <= "0101001111100100";
        wait for clk_period;
        A <= "1100011101010101";
        B <= "0010100111101111";
        C <= "0001001111111011";
        wait for clk_period;
        A <= "0001010111000101";
        B <= "1010111001110000";
        C <= "1101010101110011";
        wait for clk_period;
        A <= "0001110110111000";
        B <= "0110000100011000";
        C <= "0001101101011101";
        wait for clk_period;
        A <= "1100100001111101";
        B <= "1001101111101000";
        C <= "1100010111100001";
        wait for clk_period;
        A <= "1111010010010000";
        B <= "1100010011000010";
        C <= "0010100000111110";
        wait for clk_period;
        A <= "0100101011111000";
        B <= "1001111011101100";
        C <= "0000111011101101";
        wait for clk_period;
        A <= "0001100010001010";
        B <= "0100010001101001";
        C <= "1011000110110101";
        wait for clk_period;
        A <= "1110000000100010";
        B <= "0001101100111000";
        C <= "1110011010000110";
        wait for clk_period;
        A <= "0101101011001101";
        B <= "0000000000110000";
        C <= "0001001010100111";
        wait for clk_period;
        A <= "0100110001011101";
        B <= "0000110101101100";
        C <= "1010001000101011";
        wait for clk_period;
        A <= "1110001010101010";
        B <= "0000011011110010";
        C <= "1000000101111010";
        wait for clk_period;
        A <= "0110100100110111";
        B <= "1110000110001111";
        C <= "1111010111100101";
        wait for clk_period;
        A <= "0111000110111101";
        B <= "0001010111011000";
        C <= "1110111011011011";
        wait for clk_period;
        A <= "0100000010010001";
        B <= "0110101010110111";
        C <= "0010001110011000";
        wait for clk_period;
        A <= "0111110101011010";
        B <= "1000111010101111";
        C <= "0110000110101000";
        wait for clk_period;
        A <= "0101011010011011";
        B <= "1101111111001111";
        C <= "0110101101110110";
        wait for clk_period;
        A <= "1111110001000010";
        B <= "1101111000100010";
        C <= "1111111100101101";
        wait for clk_period;
        A <= "0000100011011011";
        B <= "1001010111001000";
        C <= "1100010111111011";
        wait for clk_period;
        A <= "0101010001001010";
        B <= "0100101001101101";
        C <= "1011011001101110";
        wait for clk_period;
        A <= "0011011101101111";
        B <= "1101110010011010";
        C <= "1000000000100111";
        wait for clk_period;
        A <= "1010100100001010";
        B <= "1111001111110110";
        C <= "1110110011011000";
        wait for clk_period;
        A <= "0010111101110100";
        B <= "1110010010010001";
        C <= "1111000011101000";
        wait for clk_period;
        A <= "1010001010001111";
        B <= "0111111101110111";
        C <= "1111000001001000";
        wait for clk_period;
        A <= "0101110110110100";
        B <= "1100001000001000";
        C <= "0110010001001010";
        wait for clk_period;
        A <= "1110000111100000";
        B <= "0111010001011011";
        C <= "0111001100110011";
        wait for clk_period;
        A <= "0001000010100010";
        B <= "0010001010110111";
        C <= "0110101000011001";
        wait for clk_period;
        A <= "0000000011101111";
        B <= "1101101010111111";
        C <= "1000000101100011";
        wait for clk_period;
        A <= "1100100111111001";
        B <= "0101000010101100";
        C <= "1011010000001010";
        wait for clk_period;
        A <= "0000010111101100";
        B <= "1010101011101101";
        C <= "1111100001010100";
        wait for clk_period;
        A <= "0010001010110001";
        B <= "1110011001010110";
        C <= "0011010111110111";
        wait for clk_period;
        A <= "0010001100111111";
        B <= "1111100101101101";
        C <= "0110111011111001";
        wait for clk_period;
        A <= "0101011001100000";
        B <= "0000011111111110";
        C <= "0010100111101010";
        wait for clk_period;
        A <= "0011000010111011";
        B <= "0011101100100101";
        C <= "1111001011010110";
        wait for clk_period;
        A <= "0100101101000111";
        B <= "0111101101001011";
        C <= "1000110001101111";
        wait for clk_period;
        A <= "0001101000001101";
        B <= "0100110011111100";
        C <= "1100011110001001";
        wait for clk_period;
        A <= "0100111101010010";
        B <= "1011100000100001";
        C <= "0111111111111101";
        wait for clk_period;
        A <= "0011010111110010";
        B <= "0010010010010010";
        C <= "0110011101110011";
        wait for clk_period;
        A <= "1011101101111100";
        B <= "1001011010011000";
        C <= "1101001001110110";
        wait for clk_period;
        A <= "0111101010111110";
        B <= "1101110111111110";
        C <= "0100010010001011";
        wait for clk_period;
        A <= "0100000000111100";
        B <= "1101011101010010";
        C <= "1100001010000011";
        wait for clk_period;
        A <= "0110101101000111";
        B <= "1001011010000000";
        C <= "1111110010101001";
        wait for clk_period;
        A <= "1111011011000001";
        B <= "1000111010000001";
        C <= "0100101010010010";
        wait for clk_period;
        A <= "1100111100010011";
        B <= "1100011111010000";
        C <= "0100110001110011";
        wait for clk_period;
        A <= "0010011101011000";
        B <= "0100001100010010";
        C <= "0111100111010111";
        wait for clk_period;
        A <= "0111011001110011";
        B <= "0101111011101101";
        C <= "0010001110000010";
        wait for clk_period;
        A <= "0100011111011101";
        B <= "0110110011110111";
        C <= "0001100011100111";
        wait for clk_period;
        A <= "0110101011111001";
        B <= "0010001001110000";
        C <= "0010010110111100";
        wait for clk_period;
        A <= "0110100011001010";
        B <= "1100001000100101";
        C <= "1111101101101111";
        wait for clk_period;
        A <= "0100111100101111";
        B <= "1111000001011111";
        C <= "0011100011011111";
        wait for clk_period;
        A <= "1000001010010010";
        B <= "0101110010001111";
        C <= "0111101001101100";
        wait for clk_period;
        A <= "1110110111101011";
        B <= "0001110000111110";
        C <= "0010101100001111";
        wait for clk_period;
        A <= "0010111010001000";
        B <= "1000001001101010";
        C <= "0110110000011001";
        wait for clk_period;
        A <= "0110111101111001";
        B <= "0110010100000111";
        C <= "0011100100001001";
        wait for clk_period;
        A <= "0000101111001000";
        B <= "1011000011100011";
        C <= "1010101010010011";
        wait for clk_period;
        A <= "1001110010110110";
        B <= "1110001010000100";
        C <= "1011110001101110";
        wait for clk_period;
        A <= "0010011001011111";
        B <= "1101011101000101";
        C <= "0101101110110011";
        wait for clk_period;
        A <= "1100100100110001";
        B <= "1110101101110011";
        C <= "1110001110011001";
        wait for clk_period;
        A <= "0011100111101101";
        B <= "0111011000010000";
        C <= "1000010011111101";
        wait for clk_period;
        A <= "1100000101011101";
        B <= "1100111001010110";
        C <= "1000010110011010";
        wait for clk_period;
        A <= "0110010010100111";
        B <= "1100010010100010";
        C <= "0111110101111110";
        wait for clk_period;
        A <= "0100001111001000";
        B <= "1001110010100111";
        C <= "1011110011001111";
        wait for clk_period;
        A <= "1100010111000011";
        B <= "0100100100100001";
        C <= "0111001001010010";
        wait for clk_period;
        A <= "0101111111011100";
        B <= "1000111001000011";
        C <= "1101001111011001";
        wait for clk_period;
        A <= "1101101001110010";
        B <= "0000000000011000";
        C <= "1110010101010101";
        wait for clk_period;
        A <= "0000101110011110";
        B <= "0111000010111011";
        C <= "1001011111000100";
        wait for clk_period;
        A <= "0110100001011110";
        B <= "1010011111100110";
        C <= "1100111001101010";
        wait for clk_period;
        A <= "0100000010111011";
        B <= "0101011010001011";
        C <= "0010101111101101";
        wait for clk_period;
        A <= "1010001101111011";
        B <= "0000000010001000";
        C <= "0101000100100000";
        wait for clk_period;
        A <= "1111000101100001";
        B <= "0101011101001011";
        C <= "1101100000100011";
        wait for clk_period;
        A <= "1101110011011101";
        B <= "0011100111101010";
        C <= "0110011101011111";
        wait for clk_period;
        A <= "0001010110011101";
        B <= "0000000101010110";
        C <= "1011101001110110";
        wait for clk_period;
        A <= "0111101100100010";
        B <= "1100110100011000";
        C <= "1101011011111100";
        wait for clk_period;
        A <= "1010111111000000";
        B <= "0010011110011101";
        C <= "1011010100100001";
        wait for clk_period;
        A <= "0010010101100000";
        B <= "0110110111010110";
        C <= "0100000100101001";
        wait for clk_period;
        A <= "1001010111010011";
        B <= "1100001110100011";
        C <= "0001101001100110";
        wait for clk_period;
        A <= "1111011000110010";
        B <= "1111101101111110";
        C <= "0000110001111011";
        wait for clk_period;
        A <= "1111100010101001";
        B <= "0100110000100100";
        C <= "0101101110110100";
        wait for clk_period;
        A <= "1101101000010001";
        B <= "0110000100100111";
        C <= "0111101000000001";
        wait for clk_period;
        A <= "1000000100001000";
        B <= "1101001101100000";
        C <= "0111100010001011";
        wait for clk_period;
        A <= "1111011100000001";
        B <= "0001011101101110";
        C <= "0111111111100000";
        wait for clk_period;
        A <= "1111010000001110";
        B <= "1010110101100001";
        C <= "1100110011010110";
        wait for clk_period;
        A <= "0100010000001101";
        B <= "0111100101111010";
        C <= "0011010111101111";
        wait for clk_period;
        A <= "1110001100000111";
        B <= "1010111100110001";
        C <= "0011110011010000";
        wait for clk_period;
        A <= "1000101010011111";
        B <= "0011010011100111";
        C <= "0101001100101111";
        wait for clk_period;
        A <= "0110000110110100";
        B <= "1010010000111110";
        C <= "0011110011100111";
        wait for clk_period;
        A <= "1111111000111100";
        B <= "0111001100101110";
        C <= "1100001101100101";
        wait for clk_period;
        A <= "1010011111110001";
        B <= "0100011100010000";
        C <= "0110101100000011";
        wait for clk_period;
        A <= "0000111111110110";
        B <= "0111111111110000";
        C <= "1011000010011111";
        wait for clk_period;
        A <= "1101010010110111";
        B <= "0100000010100001";
        C <= "0011000000000110";
        wait for clk_period;
        A <= "1110110000010010";
        B <= "1010111010000100";
        C <= "0010111111100010";
        wait for clk_period;
        A <= "0110001110111101";
        B <= "1100111001111001";
        C <= "1110000001100000";
        wait for clk_period;
        A <= "0001001111110011";
        B <= "1011010000010110";
        C <= "1010101000010001";
        wait for clk_period;
        A <= "0100101110011001";
        B <= "1111010101111111";
        C <= "1111101001110001";
        wait for clk_period;
        A <= "1100110010111010";
        B <= "0110111011101000";
        C <= "1001101111110000";
        wait for clk_period;
        A <= "0001111000011001";
        B <= "1111000001001010";
        C <= "1010111101111110";
        wait for clk_period;
        A <= "0000100111000111";
        B <= "0000111000001000";
        C <= "1001000100101001";
        wait for clk_period;
        A <= "1000110001100110";
        B <= "1101011110101100";
        C <= "1011110101011001";
        wait for clk_period;
        A <= "1000000111110010";
        B <= "1001001110101011";
        C <= "0100101101011110";
        wait for clk_period;
        A <= "0010010010011001";
        B <= "1011111110100010";
        C <= "1001010110010001";
        wait for clk_period;
        A <= "1101010000111011";
        B <= "0010010101101101";
        C <= "1010011001001101";
        wait for clk_period;
        A <= "0100100010001010";
        B <= "1001111100110111";
        C <= "0001111010111001";
        wait for clk_period;
        A <= "1100000111000101";
        B <= "1001100101110011";
        C <= "0010100010111111";
        wait for clk_period;
        A <= "1110011100110000";
        B <= "0001010011000101";
        C <= "1110001001110111";
        wait for clk_period;
        A <= "0101010010111101";
        B <= "1111101010000001";
        C <= "0101010100111101";
        wait for clk_period;
        A <= "1001011111111011";
        B <= "1110001000100110";
        C <= "1100111100001000";
        wait for clk_period;
        A <= "0011011101001000";
        B <= "1100010111001111";
        C <= "1011110100100010";
        wait for clk_period;
        A <= "0010001001011000";
        B <= "1011100111000010";
        C <= "1110100111100000";
        wait for clk_period;
        A <= "0010100101000100";
        B <= "1111010010001111";
        C <= "1110111010001011";
        wait for clk_period;
        A <= "0010110011100011";
        B <= "0110110110010010";
        C <= "1001010000010001";
        wait for clk_period;
        A <= "0110000100110100";
        B <= "0110101011011100";
        C <= "0010111111001000";
        wait for clk_period;
        A <= "1011011100000011";
        B <= "0011001011011101";
        C <= "1101111010100000";
        wait for clk_period;
        A <= "0001001110001010";
        B <= "1000100010100110";
        C <= "0001011010100111";
        wait for clk_period;
        A <= "1101011001101001";
        B <= "1010111000011100";
        C <= "1001110111100001";
        wait for clk_period;
        A <= "0110100011101111";
        B <= "1001101010100101";
        C <= "1011100001111110";
        wait for clk_period;
        A <= "1101110011111111";
        B <= "0101000011101010";
        C <= "0011100000101010";
        wait for clk_period;
        A <= "1000101110101000";
        B <= "0001100101100001";
        C <= "1101101110110011";
        wait for clk_period;
        A <= "1010101011001000";
        B <= "0100000111110101";
        C <= "1010011001110000";
        wait for clk_period;
        A <= "0101001101111100";
        B <= "1111111101101101";
        C <= "0101010011010000";
        wait for clk_period;
        A <= "0110010111000001";
        B <= "0011101000100100";
        C <= "0010111001100110";
        wait for clk_period;
        A <= "0100010110100000";
        B <= "1111011111011010";
        C <= "0000011100000110";
        wait for clk_period;
        A <= "0001001101111101";
        B <= "1010110010010010";
        C <= "1010101111110100";
        wait for clk_period;
        A <= "0110100111101100";
        B <= "1010110001000111";
        C <= "0001110110011101";
        wait for clk_period;
        A <= "0000000100101101";
        B <= "0010010011011100";
        C <= "0010110100110001";
        wait for clk_period;
        A <= "1101100011110001";
        B <= "1000110110110011";
        C <= "1000011110100101";
        wait for clk_period;
        A <= "0001111010000011";
        B <= "1001010010010010";
        C <= "1010110111011110";
        wait for clk_period;
        A <= "0101010000011101";
        B <= "1011111010010101";
        C <= "1010100001100100";
        wait for clk_period;
        A <= "1000011110011010";
        B <= "1101010110100101";
        C <= "1111010010101110";
        wait for clk_period;
        A <= "1011011111000001";
        B <= "0010111100100011";
        C <= "0110001001111000";
        wait for clk_period;
        A <= "1011110111100100";
        B <= "1100001110111001";
        C <= "0110011000011101";
        wait for clk_period;
        A <= "0001000100011001";
        B <= "0110101011110100";
        C <= "0111100100101111";
        wait for clk_period;
        A <= "1101001000010010";
        B <= "0100111000010100";
        C <= "1010011100011000";
        wait for clk_period;
        A <= "1000100000011111";
        B <= "1110010010011001";
        C <= "1101101011010011";
        wait for clk_period;
        A <= "0101111110110010";
        B <= "0111111101110101";
        C <= "1000000110000100";
        wait for clk_period;
        A <= "0011001000100001";
        B <= "1101000111010111";
        C <= "0010010101111010";
        wait for clk_period;
        A <= "0111100000101011";
        B <= "1110110011111000";
        C <= "1100100010000001";
        wait for clk_period;
        A <= "1110000110100100";
        B <= "0001100001010001";
        C <= "1111000001001101";
        wait for clk_period;
        A <= "0011011101100010";
        B <= "1001100101001100";
        C <= "1011010101110000";
        wait for clk_period;
        A <= "1010010001101000";
        B <= "1011011101100100";
        C <= "1100010001010000";
        wait for clk_period;
        A <= "1111111110011100";
        B <= "1101011010110001";
        C <= "0000100010111010";
        wait for clk_period;
        A <= "1011101010010100";
        B <= "1101100111001011";
        C <= "0000001000011100";
        wait for clk_period;
        A <= "0001010001010111";
        B <= "1100011000010110";
        C <= "0010101000001001";
        wait for clk_period;
        A <= "1110000011010110";
        B <= "0000110001111000";
        C <= "1101011110111000";
        wait for clk_period;
        A <= "1011000101010000";
        B <= "0011010111011100";
        C <= "0000010010010011";
        wait for clk_period;
        A <= "1011000111001110";
        B <= "1010101100110110";
        C <= "1101100111011001";
        wait for clk_period;
        A <= "1100011000010000";
        B <= "0000000010001011";
        C <= "0101101110111110";
        wait for clk_period;
        A <= "0000000101001011";
        B <= "0101101001110011";
        C <= "1001000000100011";
        wait for clk_period;
        A <= "0011101001011101";
        B <= "1110110011111001";
        C <= "0000000101111001";
        wait for clk_period;
        A <= "0011101111100101";
        B <= "0100011110111000";
        C <= "0110110110110101";
        wait for clk_period;
        A <= "0011101110010111";
        B <= "0010101010101010";
        C <= "0110011101111111";
        wait for clk_period;
        A <= "0001011111001001";
        B <= "0110111010010110";
        C <= "1010100110110001";
        wait for clk_period;
        A <= "1110100101110000";
        B <= "0101000100011101";
        C <= "0010110000011001";
        wait for clk_period;
        A <= "1011010100001110";
        B <= "0100111101010000";
        C <= "0100011000101001";
        wait for clk_period;
        A <= "1010101100011100";
        B <= "0001000110100111";
        C <= "0100001010110111";
        wait for clk_period;
        A <= "1010011011010110";
        B <= "0111111011111011";
        C <= "0110010101000011";
        wait for clk_period;
        A <= "0001101010110010";
        B <= "1000000100111001";
        C <= "1110000100011001";
        wait for clk_period;
        A <= "0111101101011001";
        B <= "1011000011111011";
        C <= "0110110011000010";
        wait for clk_period;
        A <= "1011101101011011";
        B <= "0100110100010100";
        C <= "0100101111111100";
        wait for clk_period;
        A <= "1000001010101001";
        B <= "0111011011110001";
        C <= "1111111100000101";
        wait for clk_period;
        A <= "0111000101010011";
        B <= "1001100000001010";
        C <= "0000100101101011";
        wait for clk_period;
        A <= "1000001000000011";
        B <= "0101100011001110";
        C <= "0101101001101110";
        wait for clk_period;
        A <= "1010101100110110";
        B <= "0111000011000000";
        C <= "0000101101110011";
        wait for clk_period;
        A <= "0111111110001010";
        B <= "0111101010111101";
        C <= "0100111010000101";
        wait for clk_period;
        A <= "1001001101001001";
        B <= "0101010011100100";
        C <= "0010110111111110";
        wait for clk_period;
        A <= "1101001010010101";
        B <= "1100100100011010";
        C <= "0010011100101011";
        wait for clk_period;
        A <= "0111100011011101";
        B <= "0010011001110110";
        C <= "1111101110100011";
        wait for clk_period;
        A <= "1010011111100010";
        B <= "1111010001011011";
        C <= "1010001010110011";
        wait for clk_period;
        A <= "0101111110000110";
        B <= "1100000000111100";
        C <= "0010110111000001";
        wait for clk_period;
        A <= "0000100100111111";
        B <= "1110001001000010";
        C <= "1110011111100000";
        wait for clk_period;
        A <= "1000001001111011";
        B <= "0101001001100000";
        C <= "1010111101011011";
        wait for clk_period;
        A <= "1000011110001011";
        B <= "1011010111011011";
        C <= "0011010110111011";
        wait for clk_period;
        A <= "1010000110001010";
        B <= "0010001111111100";
        C <= "0111000101111110";
        wait for clk_period;
        A <= "0001000101111111";
        B <= "0010010010011110";
        C <= "0000111010010100";
        wait for clk_period;
        A <= "0000110111001100";
        B <= "0100010000111001";
        C <= "0010101001010110";
        wait for clk_period;
        A <= "0011010101010000";
        B <= "0100111111110000";
        C <= "1101100101011010";
        wait for clk_period;
        A <= "1110111111010000";
        B <= "1101011010100010";
        C <= "0111101011001100";
        wait for clk_period;
        A <= "1100111001110011";
        B <= "0011101100011011";
        C <= "0101110000001010";
        wait for clk_period;
        A <= "0011100011110110";
        B <= "0101100011010011";
        C <= "1000000100100010";
        wait for clk_period;
        A <= "0001001110001110";
        B <= "1010011001111101";
        C <= "0001110111000010";
        wait for clk_period;
        A <= "1111011010000111";
        B <= "0001000011100100";
        C <= "0111111100011011";
        wait for clk_period;
        A <= "1011010011101111";
        B <= "0101000110011001";
        C <= "1000101011101110";
        wait for clk_period;
        A <= "0011010000111001";
        B <= "0001111101110111";
        C <= "1110100100001011";
        wait for clk_period;
        A <= "1001100010010000";
        B <= "1110010110010111";
        C <= "0111000110101110";
        wait for clk_period;
        A <= "1011011011101000";
        B <= "0100000100011101";
        C <= "0011101111110101";
        wait for clk_period;
        A <= "0111011110100000";
        B <= "0001101101001001";
        C <= "1001101001100001";
        wait for clk_period;
        A <= "0110011001000100";
        B <= "1110001011111010";
        C <= "1101010101000100";
        wait for clk_period;
        A <= "1100001000000001";
        B <= "1001100010000001";
        C <= "0011100010011001";
        wait for clk_period;
        A <= "1010101010001010";
        B <= "0010100001001100";
        C <= "1011011110101001";
        wait for clk_period;
        A <= "1001111000100110";
        B <= "1101000010100101";
        C <= "1010001010110100";
        wait for clk_period;
        A <= "0100011110011010";
        B <= "1010101000101100";
        C <= "1111001011010100";
        wait for clk_period;
        A <= "1011011010110010";
        B <= "1101110011010001";
        C <= "0101110010001001";
        wait for clk_period;
        A <= "0011011111100101";
        B <= "1010101110100011";
        C <= "1010111000000100";
        wait for clk_period;
        A <= "1010111100001001";
        B <= "0110001010110011";
        C <= "1001010011100010";
        wait for clk_period;
        A <= "0001100011011000";
        B <= "0000101110011000";
        C <= "0101010100001000";
        wait for clk_period;
        A <= "0001110100110011";
        B <= "0101100110111001";
        C <= "1010100100111001";
        wait for clk_period;
        A <= "1100111101001101";
        B <= "1001101111110101";
        C <= "0100001101010011";
        wait for clk_period;
        A <= "1001011110111011";
        B <= "0111011001101010";
        C <= "0010000101110111";
        wait for clk_period;
        A <= "1101101000101000";
        B <= "0100010111000110";
        C <= "0100000000111100";
        wait for clk_period;
        A <= "1011001001011000";
        B <= "1111110111101100";
        C <= "1011111111100111";
        wait for clk_period;
        A <= "1011001110000011";
        B <= "0101110100010100";
        C <= "1000010000111010";
        wait for clk_period;
        A <= "1011010111010100";
        B <= "1011011100100110";
        C <= "0101000101111101";
        wait for clk_period;
        A <= "1110000011101110";
        B <= "0111011000000001";
        C <= "0000100110110110";
        wait for clk_period;
        A <= "0000011011001100";
        B <= "1111001110001010";
        C <= "1100000001001110";
        wait for clk_period;
        A <= "1110111000110110";
        B <= "1110101111001100";
        C <= "1101110010100010";
        wait for clk_period;
        A <= "1000000000110110";
        B <= "1111111011100111";
        C <= "1100111100111101";
        wait for clk_period;
        A <= "1000001010000111";
        B <= "1111111010111000";
        C <= "1100111010010100";
        wait for clk_period;
        A <= "1100100101011011";
        B <= "1011010010000000";
        C <= "1101101100011110";
        wait for clk_period;
        A <= "1010011110000110";
        B <= "1101111100111010";
        C <= "0000001111000101";
        wait for clk_period;
        A <= "0010011010001011";
        B <= "1101110110000111";
        C <= "1100011100011000";
        wait for clk_period;
        A <= "1010111011110000";
        B <= "1100001000110110";
        C <= "1000110001101101";
        wait for clk_period;
        A <= "1011110010011001";
        B <= "1001011100001000";
        C <= "1011000010000001";
        wait for clk_period;
        A <= "1000011110001011";
        B <= "0010001101000100";
        C <= "0010001100110000";
        wait for clk_period;
        A <= "0100100010010011";
        B <= "1110100100110100";
        C <= "0010100010110011";
        wait for clk_period;
        A <= "1000110101101000";
        B <= "1100110101100000";
        C <= "1100000001100000";
        wait for clk_period;
        A <= "1110011001000001";
        B <= "1011110010001101";
        C <= "1000011010101011";
        wait for clk_period;
        A <= "1111000100111101";
        B <= "1110011011101001";
        C <= "1111100111101110";
        wait for clk_period;
        A <= "0100010100000000";
        B <= "0010010010110101";
        C <= "0011000011101001";
        wait for clk_period;
        A <= "1001010111101111";
        B <= "1000100000000010";
        C <= "0101111111101001";
        wait for clk_period;
        A <= "1110010100111000";
        B <= "0011011010101010";
        C <= "0001000001000001";
        wait for clk_period;
        A <= "0111000100001100";
        B <= "0001101000001101";
        C <= "1000000011110100";
        wait for clk_period;
        A <= "0111001101110110";
        B <= "0111111110010101";
        C <= "1100101001011101";
        wait for clk_period;
        A <= "1110111000100010";
        B <= "0011011000101000";
        C <= "1010000000110100";
        wait for clk_period;
        A <= "1111111001010000";
        B <= "1100011010110111";
        C <= "1111100111000010";
        wait for clk_period;
        A <= "0010010100110110";
        B <= "0000010000110110";
        C <= "0110110000110011";
        wait for clk_period;
        A <= "0001010100111001";
        B <= "1000100101110110";
        C <= "1101011110101111";
        wait for clk_period;
        A <= "1101101111111110";
        B <= "1110001100111011";
        C <= "0001110001100001";
        wait for clk_period;
        A <= "0100000110110011";
        B <= "1110011111010111";
        C <= "0000001001100100";
        wait for clk_period;
        A <= "1000000111101011";
        B <= "0011111111010100";
        C <= "0011110000010111";
        wait for clk_period;
        A <= "1000101111101110";
        B <= "1001001110000101";
        C <= "0001011000100000";
        wait for clk_period;
        A <= "1001111000100101";
        B <= "0101101101011011";
        C <= "1000111111111111";
        wait for clk_period;
        A <= "1111101010000101";
        B <= "0100000110110011";
        C <= "0001001111111010";
        wait for clk_period;
        A <= "1000000111010011";
        B <= "1100101100010011";
        C <= "1010010000110100";
        wait for clk_period;
        A <= "0010100010010101";
        B <= "0111000001001101";
        C <= "1111100111110010";
        wait for clk_period;
        A <= "1100001111101011";
        B <= "1000100001011111";
        C <= "0011101011110000";
        wait for clk_period;
        A <= "0000010100110111";
        B <= "0010010100010001";
        C <= "0111100011100011";
        wait for clk_period;
        A <= "0101010001010110";
        B <= "0001011101100101";
        C <= "0001111011100001";
        wait for clk_period;
        A <= "1101101101010111";
        B <= "0000110011100110";
        C <= "1111111000100000";
        wait for clk_period;
        A <= "1010011101100110";
        B <= "1001101111100000";
        C <= "1001111001010011";
        wait for clk_period;
        A <= "0001110111100000";
        B <= "0000000000010100";
        C <= "0001100111011110";
        wait for clk_period;
        A <= "1010000000101100";
        B <= "1010001010100101";
        C <= "1111011001010111";
        wait for clk_period;
        A <= "0010101100001100";
        B <= "1110001110101010";
        C <= "0000101000100000";
        wait for clk_period;
        A <= "1000111110011101";
        B <= "1001111010011011";
        C <= "1100010011010000";
        wait for clk_period;
        A <= "0001101001111011";
        B <= "0011110111101100";
        C <= "1101110011001101";
        wait for clk_period;
        A <= "1100101110111001";
        B <= "0100010100010111";
        C <= "0101010110100100";
        wait for clk_period;
        A <= "1111101110101111";
        B <= "0011111011000100";
        C <= "1101000000001101";
        wait for clk_period;
        A <= "1010110010011000";
        B <= "0010100111101100";
        C <= "0111101001001001";
        wait for clk_period;
        A <= "0100111110100101";
        B <= "1000111011011011";
        C <= "1011101010110011";
        wait for clk_period;
        A <= "1000111010111000";
        B <= "1000010111010100";
        C <= "0010010111100010";
        wait for clk_period;
        A <= "1010101101100010";
        B <= "1101111010001000";
        C <= "0101001111001100";
        wait for clk_period;
        A <= "0111001111000001";
        B <= "1001010100011101";
        C <= "0110001100011011";
        wait for clk_period;
        A <= "1011000111101101";
        B <= "0100001011000100";
        C <= "0010010011001001";
        wait for clk_period;
        A <= "0011000001001011";
        B <= "0110111111100000";
        C <= "1011000110110011";
        wait for clk_period;
        A <= "1111101110001011";
        B <= "1110110111101001";
        C <= "0110000011110000";
        wait for clk_period;
        A <= "0110010011010111";
        B <= "0111111000110100";
        C <= "1110101001100010";
        wait for clk_period;
        A <= "1110001111000010";
        B <= "0000000000100111";
        C <= "0110100010100110";
        wait for clk_period;
        A <= "1010101000001111";
        B <= "1100110011101100";
        C <= "0000100011001101";
        wait for clk_period;
        A <= "0001111000101011";
        B <= "0010000001101011";
        C <= "0010001010110100";
        wait for clk_period;
        A <= "0111110010101011";
        B <= "1110100001100101";
        C <= "0110101010000100";
        wait for clk_period;
        A <= "0111110010100011";
        B <= "0100110010010111";
        C <= "0010000100101001";
        wait for clk_period;
        A <= "0111110101011011";
        B <= "1001010001101000";
        C <= "1010110010010100";
        wait for clk_period;
        A <= "1101100110111110";
        B <= "0000101011000111";
        C <= "1101011100010000";
        wait for clk_period;
        A <= "1000000000001101";
        B <= "1011111010111110";
        C <= "1000110100110111";
        wait for clk_period;
        A <= "1100001110000100";
        B <= "0101100111001110";
        C <= "0000011010011010";
        wait for clk_period;
        A <= "1101001000010001";
        B <= "1100000101001000";
        C <= "1111101100100011";
        wait for clk_period;
        A <= "0000010010100111";
        B <= "1110111110000011";
        C <= "1110001001111110";
        wait for clk_period;
        A <= "0011001110010110";
        B <= "0010110101101100";
        C <= "0110000110010000";
        wait for clk_period;
        A <= "1010010010110000";
        B <= "0110011110100111";
        C <= "1101101110111110";
        wait for clk_period;
        A <= "1011100100110100";
        B <= "0001010110000111";
        C <= "0110110010110101";
        wait for clk_period;
        A <= "0011010100111010";
        B <= "0011001110011011";
        C <= "1110011011001001";
        wait for clk_period;
        A <= "0011100010100110";
        B <= "0110000001101010";
        C <= "0011101100011111";
        wait for clk_period;
        A <= "1010010001110000";
        B <= "1111100000000110";
        C <= "1000101000000101";
        wait for clk_period;
        A <= "1000001101111000";
        B <= "1010111110001110";
        C <= "1101100110110000";
        wait for clk_period;
        A <= "1000010100101010";
        B <= "0001101110010011";
        C <= "1000101111101011";
        wait for clk_period;
        A <= "1111000010011001";
        B <= "1011100110111011";
        C <= "1111001010101011";
        wait for clk_period;
        A <= "0011111100101010";
        B <= "1101000011100111";
        C <= "0100100110110011";
        wait for clk_period;
        A <= "0111011001000101";
        B <= "1000111010101011";
        C <= "1001010000110110";
        wait for clk_period;
        A <= "1100101010110100";
        B <= "0001000100101000";
        C <= "0101011001000100";
        wait for clk_period;
        A <= "1011000011000000";
        B <= "0011011100010110";
        C <= "0010000000100000";
        wait for clk_period;
        A <= "0101010010001010";
        B <= "0010010011100001";
        C <= "1000101000000001";
        wait for clk_period;
        A <= "1010011110100110";
        B <= "0001111111001111";
        C <= "1100110100001110";
        wait for clk_period;
        A <= "0110000110111001";
        B <= "0010011000111101";
        C <= "0111111011101010";
        wait for clk_period;
        A <= "0011110010001111";
        B <= "1001111000000100";
        C <= "1100011100101001";
        wait for clk_period;
        A <= "0010100110001110";
        B <= "0111101011000100";
        C <= "1000100101110010";
        wait for clk_period;
        A <= "1001011110101100";
        B <= "0001100010110100";
        C <= "0100110111100010";
        wait for clk_period;
        A <= "1111100000001010";
        B <= "0100111000000101";
        C <= "1011011100000001";
        wait for clk_period;
        A <= "1001001101010010";
        B <= "0001001010011110";
        C <= "1010001110111111";
        wait for clk_period;
        A <= "1000111000010111";
        B <= "0111110011110101";
        C <= "1001111100110101";
        wait for clk_period;
        A <= "1001111100110000";
        B <= "1110101101101111";
        C <= "0111100100001011";
        wait for clk_period;
        A <= "1000110000010100";
        B <= "1110011001101100";
        C <= "1010011010001001";
        wait for clk_period;
        A <= "1010000000000100";
        B <= "1000100011100100";
        C <= "0101010001111000";
        wait for clk_period;
        A <= "1100001111111100";
        B <= "1101110010011111";
        C <= "1011010110010001";
        wait for clk_period;
        A <= "1100010011010001";
        B <= "0011010101111011";
        C <= "0100000010100011";
        wait for clk_period;
        A <= "1101110110101010";
        B <= "0001011100111000";
        C <= "0110010010100111";
        wait for clk_period;
        A <= "1011000100000010";
        B <= "0101000101111011";
        C <= "1111111101001000";
        wait for clk_period;
        A <= "0011000000001011";
        B <= "1000010100000000";
        C <= "1011110100001110";
        wait for clk_period;
        A <= "0100000000110111";
        B <= "1100000011101011";
        C <= "1001001110011000";
        wait for clk_period;
        A <= "1011100011100000";
        B <= "0010001111100111";
        C <= "0101100111110111";
        wait for clk_period;
        A <= "1101010010100111";
        B <= "0101111001101010";
        C <= "0000111100001110";
        wait for clk_period;
        A <= "0001110111000110";
        B <= "0101101111001100";
        C <= "0110001011001010";
        wait for clk_period;
        A <= "1110001111001100";
        B <= "0000011010010000";
        C <= "1101001001000001";
        wait for clk_period;
        A <= "0100100010000010";
        B <= "0111000000001100";
        C <= "0100001101110011";
        wait for clk_period;
        A <= "0000110110111011";
        B <= "0110000010010000";
        C <= "1001111011100111";
        wait for clk_period;
        A <= "0011011011011010";
        B <= "0101010011110111";
        C <= "1101101111111111";
        wait for clk_period;
        A <= "0011011101000110";
        B <= "1000100001010100";
        C <= "0110000110011101";
        wait for clk_period;
        A <= "0110000010001010";
        B <= "0101101000110101";
        C <= "0000010101111010";
        wait for clk_period;
        A <= "0101001100111111";
        B <= "0111111000000100";
        C <= "0100100001001111";
        wait for clk_period;
        A <= "1011011001101101";
        B <= "0010110101010111";
        C <= "0100101001110011";
        wait for clk_period;
        A <= "0000110000010100";
        B <= "0010011000111011";
        C <= "1000001010110011";
        wait for clk_period;
        A <= "0011000001000000";
        B <= "1100110100110010";
        C <= "0001010011001001";
        wait for clk_period;
        A <= "0011100110100111";
        B <= "1101000101010111";
        C <= "0010110001111011";
        wait for clk_period;
        A <= "0101101001000101";
        B <= "0100110010010010";
        C <= "0110010011001010";
        wait for clk_period;
        A <= "1011100110000110";
        B <= "0101011010101010";
        C <= "0000101100100101";
        wait for clk_period;
        A <= "0100101111100011";
        B <= "1101010101000010";
        C <= "1100011001100000";
        wait for clk_period;
        A <= "1110001001111111";
        B <= "1100001011001111";
        C <= "0010001001100101";
        wait for clk_period;
        A <= "1001001011000010";
        B <= "0000001010110011";
        C <= "1011111101011101";
        wait for clk_period;
        A <= "0000101011011011";
        B <= "0011001011011000";
        C <= "1011101100110110";
        wait for clk_period;
        A <= "1010101111110100";
        B <= "1010100011000100";
        C <= "0100000000111011";
        wait for clk_period;
        A <= "0101001110110011";
        B <= "1011100110111010";
        C <= "1110010000110011";
        wait for clk_period;
        A <= "0010111110000110";
        B <= "0010000101011011";
        C <= "0100111011001010";
        wait for clk_period;
        A <= "0000010011110111";
        B <= "0110110011110111";
        C <= "1110011100011001";
        wait for clk_period;
        A <= "1011110000101001";
        B <= "0000001110110110";
        C <= "1111110111101101";
        wait for clk_period;
        A <= "1000111000001111";
        B <= "1011010010111011";
        C <= "1010011000011101";
        wait for clk_period;
        A <= "0100000000010111";
        B <= "1111100011000111";
        C <= "0011001111000001";
        wait for clk_period;
        A <= "1011100100110010";
        B <= "1011011110000010";
        C <= "0010100100111010";
        wait for clk_period;
        A <= "0100101110100101";
        B <= "1010011110010000";
        C <= "0100001011111101";
        wait for clk_period;
        A <= "0100011111111001";
        B <= "1111001000011001";
        C <= "1001101000011000";
        wait for clk_period;
        A <= "0001001010011011";
        B <= "1101010111010001";
        C <= "0010001010011011";
        wait for clk_period;
        A <= "0110110111001110";
        B <= "0100111100110100";
        C <= "0111100111101010";
        wait for clk_period;
        A <= "0110101010100010";
        B <= "1001010001101101";
        C <= "0101000000110010";
        wait for clk_period;
        A <= "0100101111100011";
        B <= "1111111011111010";
        C <= "1101111100101111";
        wait for clk_period;
        A <= "1000101101000000";
        B <= "1111000101000000";
        C <= "0011011100011000";
        wait for clk_period;
        A <= "0101011111001011";
        B <= "0111111110001101";
        C <= "0011101010000101";
        wait for clk_period;
        A <= "1100011010110111";
        B <= "0011000101111111";
        C <= "1010110010100101";
        wait for clk_period;
        A <= "0001001010000111";
        B <= "1010011101111100";
        C <= "1111011110100000";
        wait for clk_period;
        A <= "1101001100011101";
        B <= "0111000110100001";
        C <= "1001100110011111";
        wait for clk_period;
        A <= "0110111011000111";
        B <= "0100110011110001";
        C <= "0000011100010000";
        wait for clk_period;
        A <= "0010001010110110";
        B <= "0111010101101000";
        C <= "0111100000111111";
        wait for clk_period;
        A <= "0110110010100001";
        B <= "1101111101000111";
        C <= "0000100100000110";
        wait for clk_period;
        A <= "1110010111101000";
        B <= "0111010001000011";
        C <= "0010011011110011";
        wait for clk_period;
        A <= "1010110101110110";
        B <= "1101010111111111";
        C <= "1101110010111001";
        wait for clk_period;
        A <= "1001101000110110";
        B <= "1111010100100011";
        C <= "1110001011010000";
        wait for clk_period;
        A <= "1111000001000000";
        B <= "1010011111000110";
        C <= "0111001011000111";
        wait for clk_period;
        A <= "0111001110011110";
        B <= "0010011001100110";
        C <= "0101111010111010";
        wait for clk_period;
        A <= "1011001001101110";
        B <= "0100101110000010";
        C <= "0010101110000001";
        wait for clk_period;
        A <= "1000010010000110";
        B <= "1110000110011001";
        C <= "0001000001110100";
        wait for clk_period;
        A <= "1011010000011010";
        B <= "0011001010001001";
        C <= "1110100101101000";
        wait for clk_period;
        A <= "0000000001111101";
        B <= "1011100001010001";
        C <= "1001101000101010";
        wait for clk_period;
        A <= "0011110111111010";
        B <= "1001010010111001";
        C <= "0100101010100000";
        wait for clk_period;
        A <= "0111111010001111";
        B <= "1101111000001111";
        C <= "0110001100000100";
        wait for clk_period;
        A <= "1010101011000000";
        B <= "1110100111010111";
        C <= "0101011010111001";
        wait for clk_period;
        A <= "1000011000000100";
        B <= "1010010010011110";
        C <= "0111011101111111";
        wait for clk_period;
        A <= "0000001101001010";
        B <= "0011011100001111";
        C <= "0101010111100010";
        wait for clk_period;
        A <= "0100100010110101";
        B <= "0000011101001011";
        C <= "0110111111111111";
        wait for clk_period;
        A <= "1100010101101011";
        B <= "1001010111000011";
        C <= "1010010000011110";
        wait for clk_period;
        A <= "1101010001001110";
        B <= "0001110110100111";
        C <= "1110100111110001";
        wait for clk_period;
        A <= "1011001001111100";
        B <= "1111010100101010";
        C <= "1111110010000010";
        wait for clk_period;
        A <= "0010111101100011";
        B <= "1110001010110001";
        C <= "1101000100100101";
        wait for clk_period;
        A <= "1011111000001001";
        B <= "0111011000000101";
        C <= "0011001100000000";
        wait for clk_period;
        A <= "0010010101110010";
        B <= "0011100001110101";
        C <= "1111101110011110";
        wait for clk_period;
        A <= "0000010001000101";
        B <= "1110101011011000";
        C <= "1110010100000000";
        wait for clk_period;
        A <= "1101010111111110";
        B <= "0111100111111000";
        C <= "0000011100111000";
        wait for clk_period;
        A <= "0101010001100111";
        B <= "0001011110010100";
        C <= "1110111000100111";
        wait for clk_period;
        A <= "0001001011110110";
        B <= "1001001111110001";
        C <= "0100100111001100";
        wait for clk_period;
        A <= "1110101001111111";
        B <= "1110110110111010";
        C <= "0010101110000011";
        wait for clk_period;
        A <= "1000100111001011";
        B <= "0101110001000000";
        C <= "1110111110001011";
        wait for clk_period;
        A <= "1010000111110101";
        B <= "1111110011100001";
        C <= "1001110100001010";
        wait for clk_period;
        A <= "0001001101000000";
        B <= "1101101110011110";
        C <= "0001001001100111";
        wait for clk_period;
        A <= "1000111100011111";
        B <= "1000100011111111";
        C <= "0101111111101110";
        wait for clk_period;
        A <= "0101001010001101";
        B <= "1000000110100011";
        C <= "1110010100111000";
        wait for clk_period;
        A <= "0000011011101110";
        B <= "0000011101111010";
        C <= "0011011010110101";
        wait for clk_period;
        A <= "0111100101111101";
        B <= "0100101010110101";
        C <= "0111001100110000";
        wait for clk_period;
        A <= "1110011111011110";
        B <= "1101000001010001";
        C <= "1101110100001000";
        wait for clk_period;
        A <= "1101110011111110";
        B <= "1011111111000010";
        C <= "1000011010100010";
        wait for clk_period;
        A <= "1100101110110101";
        B <= "0111100110000100";
        C <= "0100000111100011";
        wait for clk_period;
        A <= "1001100000000011";
        B <= "0111100110100101";
        C <= "1111111011001001";
        wait for clk_period;
        A <= "1101000011010011";
        B <= "0100110111100011";
        C <= "0011101100100010";
        wait for clk_period;
        A <= "1000010010010001";
        B <= "0101000001110011";
        C <= "1110101101001011";
        wait for clk_period;
        A <= "0010000001111111";
        B <= "1001110110101011";
        C <= "0011101111100111";
        wait for clk_period;
        A <= "0001101100010101";
        B <= "0101000110111111";
        C <= "0110101100110001";
        wait for clk_period;
        A <= "0001100000100110";
        B <= "1100011001110011";
        C <= "1111101111100101";
        wait for clk_period;
        A <= "0110111110110001";
        B <= "0111110111111011";
        C <= "0001010111011011";
        wait for clk_period;
        A <= "0011101100010101";
        B <= "0011110001011100";
        C <= "1110000111110111";
        wait for clk_period;
        A <= "0101011100011101";
        B <= "1010000100101010";
        C <= "1100110010000111";
        wait for clk_period;
        A <= "1000011100000010";
        B <= "0101100110011010";
        C <= "1011110001111100";
        wait for clk_period;
        A <= "1011011000001011";
        B <= "1110101100010000";
        C <= "1010001010110111";
        wait for clk_period;
        A <= "0101000100110100";
        B <= "0101001101101100";
        C <= "0000100111100100";
        wait for clk_period;
        A <= "1011101011110010";
        B <= "0100001100100001";
        C <= "0110111100010110";
        wait for clk_period;
        A <= "1110000100011011";
        B <= "0110000000110011";
        C <= "0010011000110111";
        wait for clk_period;
        A <= "1011100010111011";
        B <= "0101111100001010";
        C <= "0001000101111100";
        wait for clk_period;
        A <= "0000001010011000";
        B <= "1101101111100111";
        C <= "1111111110011100";
        wait for clk_period;
        A <= "0001000010011111";
        B <= "1110110011110000";
        C <= "0010001010111010";
        wait for clk_period;
        A <= "0110111101011010";
        B <= "1111010001010111";
        C <= "0011000001101001";
        wait for clk_period;
        A <= "1110100011011111";
        B <= "0111101111111100";
        C <= "1101011101110001";
        wait for clk_period;
        A <= "0001101000010001";
        B <= "1000010010110000";
        C <= "1111101010011110";
        wait for clk_period;
        A <= "1100101111100101";
        B <= "0110000110011110";
        C <= "1110010100010011";
        wait for clk_period;
        A <= "0101011101110101";
        B <= "0010000110001111";
        C <= "1100111010011111";
        wait for clk_period;
        A <= "1010100111000101";
        B <= "1010000000101011";
        C <= "0011110010100100";
        wait for clk_period;
        A <= "0101100101100010";
        B <= "0101111011011011";
        C <= "1111010010000001";
        wait for clk_period;
        A <= "1000101100111100";
        B <= "1100111011000010";
        C <= "1110111001110110";
        wait for clk_period;
        A <= "1111101111001110";
        B <= "0010001010000101";
        C <= "0101110101011101";
        wait for clk_period;
        A <= "0010111110010010";
        B <= "0101100101111011";
        C <= "0101000101101100";
        wait for clk_period;
        A <= "1111010100110010";
        B <= "1101010011010111";
        C <= "0000110000110100";
        wait for clk_period;
        A <= "0010010101010011";
        B <= "0011101110000101";
        C <= "0111011000111100";
        wait for clk_period;
        A <= "0011011110001110";
        B <= "0011000000010000";
        C <= "1110110111011011";
        wait for clk_period;
        A <= "1110101011000100";
        B <= "1001011010011011";
        C <= "1001111101101001";
        wait for clk_period;
        A <= "0011011110100110";
        B <= "1011011101101000";
        C <= "0111000000001001";
        wait for clk_period;
        A <= "0000110100101101";
        B <= "1011100101100101";
        C <= "1010111101000001";
        wait for clk_period;
        A <= "0011110110000011";
        B <= "1101110001101111";
        C <= "0001011111110100";
        wait for clk_period;
        A <= "1111000000111100";
        B <= "0110111010010010";
        C <= "0101001011000100";
        wait for clk_period;
        A <= "0000010011011101";
        B <= "1011100011100100";
        C <= "1111000010111111";
        wait for clk_period;
        A <= "1010001011010011";
        B <= "0111010111100010";
        C <= "1001010001011001";
        wait for clk_period;
        A <= "0100001110010010";
        B <= "0000110101101100";
        C <= "1001100110100111";
        wait for clk_period;
        A <= "0011011110110000";
        B <= "1100101110011010";
        C <= "0011100110000001";
        wait for clk_period;
        A <= "0111101100001011";
        B <= "0011010011101010";
        C <= "0100101000001001";
        wait for clk_period;
        A <= "1100001001011001";
        B <= "0111110111000001";
        C <= "1111111010010111";
        wait for clk_period;
        A <= "1111010111111000";
        B <= "0010111001101001";
        C <= "1010110100111010";
        wait for clk_period;
        A <= "1110011011010110";
        B <= "0101010111011101";
        C <= "1101011000000110";
        wait for clk_period;
        A <= "0100011010001001";
        B <= "1100111100110100";
        C <= "0001110010010110";
        wait for clk_period;
        A <= "1110110101011001";
        B <= "0101111101010111";
        C <= "0111111000010010";
        wait for clk_period;
        A <= "0010010000000010";
        B <= "1101010011010111";
        C <= "0001101100101101";
        wait for clk_period;
        A <= "1101100000010111";
        B <= "0001001001000001";
        C <= "0011011100001010";
        wait for clk_period;
        A <= "0001011110100000";
        B <= "1100110111101000";
        C <= "1000001001011010";
        wait for clk_period;
        A <= "1010110001100110";
        B <= "0001011001101101";
        C <= "0000001011010001";
        wait for clk_period;
        A <= "0011101001000111";
        B <= "1010011110101100";
        C <= "1011100100011001";
        wait for clk_period;
        A <= "0001011011010100";
        B <= "1010111010000010";
        C <= "0011011101100111";
        wait for clk_period;
        A <= "1100011100111000";
        B <= "0010010011111110";
        C <= "0111101100111010";
        wait for clk_period;
        A <= "1111100001010010";
        B <= "0110010010110111";
        C <= "0011100101011010";
        wait for clk_period;
        A <= "1000110010000111";
        B <= "1000001110000111";
        C <= "1100110001010000";
        wait for clk_period;
        A <= "1000100101010101";
        B <= "0000110111000100";
        C <= "1010001010110001";
        wait for clk_period;
        A <= "0110111001010011";
        B <= "0001001111100110";
        C <= "1000101010101011";
        wait for clk_period;
        A <= "1001000011000000";
        B <= "1001100101001001";
        C <= "0010011000001011";
        wait for clk_period;
        A <= "1100100001100111";
        B <= "0101110011011011";
        C <= "1000000101110010";
        wait for clk_period;
        A <= "0110010101001001";
        B <= "0101111110100011";
        C <= "0001111001011000";
        wait for clk_period;
        A <= "1000010000111000";
        B <= "1110101001011011";
        C <= "1000101011001111";
        wait for clk_period;
        A <= "0110010110111001";
        B <= "1000101100101010";
        C <= "0000010000011111";
        wait for clk_period;
        A <= "0100100000011100";
        B <= "0101000110000100";
        C <= "1111011100011001";
        wait for clk_period;
        A <= "1101010010010010";
        B <= "0100010010101000";
        C <= "1101010000011111";
        wait for clk_period;
        A <= "1100001101001110";
        B <= "1010001000000111";
        C <= "1101110111000001";
        wait for clk_period;
        A <= "0010010011101001";
        B <= "0111000010100101";
        C <= "1010011101010110";
        wait for clk_period;
        A <= "1111110101111101";
        B <= "0011110111010001";
        C <= "1111000000100100";
        wait for clk_period;
        A <= "1101011110011110";
        B <= "0111001111101010";
        C <= "0011111000011110";
        wait for clk_period;
        A <= "1000001000110010";
        B <= "0110000101000001";
        C <= "0000001000000011";
        wait for clk_period;
        A <= "1011001101010010";
        B <= "0010000001111011";
        C <= "0100100010110001";
        wait for clk_period;
        A <= "1111011110111100";
        B <= "1111110001111101";
        C <= "0000111000010001";
        wait for clk_period;
        A <= "1110001000100101";
        B <= "0000010101001001";
        C <= "0100111101110010";
        wait for clk_period;
        A <= "1011001101011011";
        B <= "0100010111001011";
        C <= "1011010101000110";
        wait for clk_period;
        A <= "0010111010100010";
        B <= "0111111010011111";
        C <= "1110001110000110";
        wait for clk_period;
        A <= "1111110110101001";
        B <= "1000011110010011";
        C <= "0000011100011000";
        wait for clk_period;
        A <= "0110110111111111";
        B <= "0101110000110000";
        C <= "0110010110110001";
        wait for clk_period;
        A <= "0100110110100000";
        B <= "1111000111100111";
        C <= "0010111110010111";
        wait for clk_period;
        A <= "0101100101110110";
        B <= "1111100011001010";
        C <= "1111111000001000";
        wait for clk_period;
        A <= "0010001101110101";
        B <= "1101101110001111";
        C <= "1100110101011010";
        wait for clk_period;
        A <= "0111011111001100";
        B <= "1011110001000100";
        C <= "0011001000101010";
        wait for clk_period;
        A <= "0011110010000101";
        B <= "1100111010100111";
        C <= "1101000001100110";
        wait for clk_period;
        A <= "1110110010101101";
        B <= "0111110010100100";
        C <= "1000010111001101";
        wait for clk_period;
        A <= "0100111100101000";
        B <= "0111001000110001";
        C <= "1001110001100001";
        wait for clk_period;
        A <= "1000110101100011";
        B <= "1100111011111110";
        C <= "1010000110010011";
        wait for clk_period;
        A <= "0101100111111010";
        B <= "1000011000010111";
        C <= "1111001010001111";
        wait for clk_period;
        A <= "1001001100111010";
        B <= "1000011000110000";
        C <= "0100011011111011";
        wait for clk_period;
        A <= "0001001011000110";
        B <= "0101010001011100";
        C <= "0101101001000110";
        wait for clk_period;
        A <= "1101101001101001";
        B <= "0011001010111101";
        C <= "0101011001001000";
        wait for clk_period;
        A <= "1000000111100011";
        B <= "0101000110000100";
        C <= "1010100001111001";
        wait for clk_period;
        A <= "0111000101011100";
        B <= "0001000000001010";
        C <= "0000001001010010";
        wait for clk_period;
        A <= "0000100011100100";
        B <= "1010101010001101";
        C <= "1110100101010011";
        wait for clk_period;
        A <= "1110000001011001";
        B <= "1001010100010101";
        C <= "0100001100011100";
        wait for clk_period;
        A <= "0000010011010110";
        B <= "1001010010000001";
        C <= "1010000100100001";
        wait for clk_period;
        A <= "0001110101001111";
        B <= "1000101110110100";
        C <= "0010111101000011";
        wait for clk_period;
        A <= "0101111010001001";
        B <= "1010100011000011";
        C <= "1001101010110100";
        wait for clk_period;
        A <= "0111010100001011";
        B <= "1111111111000111";
        C <= "1101100011010000";
        wait for clk_period;
        A <= "0100000010001100";
        B <= "0111011000000000";
        C <= "0010111011010000";
        wait for clk_period;
        A <= "0000000110101001";
        B <= "0100001100111011";
        C <= "0011110100101001";
        wait for clk_period;
        A <= "1001110010011011";
        B <= "0111011001111100";
        C <= "1000100010010000";
        wait for clk_period;
        A <= "1101101101001001";
        B <= "0100011101111001";
        C <= "1011111110111110";
        wait for clk_period;
        A <= "0010100101001110";
        B <= "1101000111011101";
        C <= "0001000101011001";
        wait for clk_period;
        A <= "0011010010110111";
        B <= "1011111100111011";
        C <= "1010010001001011";
        wait for clk_period;
        A <= "0101100000001110";
        B <= "1010101101000110";
        C <= "1101010111010110";
        wait for clk_period;
        A <= "0100000010101001";
        B <= "0011100100001011";
        C <= "1100100100011100";
        wait for clk_period;
        A <= "0111111110010110";
        B <= "0111100011111101";
        C <= "1110000010110011";
        wait for clk_period;
        A <= "0101011011001110";
        B <= "1111101100110010";
        C <= "0100010010100001";
        wait for clk_period;
        A <= "1000011011101100";
        B <= "0110100110101010";
        C <= "0111010001001101";
        wait for clk_period;
        A <= "0111110100010011";
        B <= "1000101001100101";
        C <= "0011100011000110";
        wait for clk_period;
        A <= "0110000110101001";
        B <= "0110001011010011";
        C <= "1011100000011000";
        wait for clk_period;
        A <= "0111111011000000";
        B <= "1010001111011011";
        C <= "0100111011100011";
        wait for clk_period;
        A <= "1011000111110000";
        B <= "1111110100100110";
        C <= "0000100001000110";
        wait for clk_period;
        A <= "0000000011001001";
        B <= "1110011101110011";
        C <= "0101000110100110";
        wait for clk_period;
        A <= "0111011111011000";
        B <= "1111101100000001";
        C <= "0011011111111110";
        wait for clk_period;
        A <= "1100110010000111";
        B <= "0110010000101111";
        C <= "1111000111111001";
        wait for clk_period;
        A <= "1111000100101000";
        B <= "0000101001000001";
        C <= "0110101010001000";
        wait for clk_period;
        A <= "0011110100000101";
        B <= "1011111110111010";
        C <= "0110001001010000";
        wait for clk_period;
        A <= "0001001100000010";
        B <= "1101011100111110";
        C <= "1000100100010011";
        wait for clk_period;
        A <= "0100100010101000";
        B <= "0100101100100111";
        C <= "0110101010101000";
        wait for clk_period;
        A <= "0000011001100111";
        B <= "0001111101100001";
        C <= "0110101000011000";
        wait for clk_period;
        A <= "1011101011010110";
        B <= "1110111010101000";
        C <= "0011101001101011";
        wait for clk_period;
        A <= "1000100110001111";
        B <= "1100101110010111";
        C <= "1011000001101001";
        wait for clk_period;
        A <= "1101111010101000";
        B <= "1010010011000101";
        C <= "1011010011010011";
        wait for clk_period;
        A <= "1111000101111011";
        B <= "1100110111000011";
        C <= "1100001100001001";
        wait for clk_period;
        A <= "1101010010100011";
        B <= "1011010111111110";
        C <= "0011101100101000";
        wait for clk_period;
        A <= "1111010101111111";
        B <= "1111010000101110";
        C <= "0010011101101101";
        wait for clk_period;
        A <= "1111011010101111";
        B <= "1100001100100000";
        C <= "0011010111011110";
        wait for clk_period;
        A <= "1011011011100101";
        B <= "0111101001101010";
        C <= "0001010100000101";
        wait for clk_period;
        A <= "1000110001111001";
        B <= "1011101111011011";
        C <= "0001001111000111";
        wait for clk_period;
        A <= "0110100011101000";
        B <= "0110100101111111";
        C <= "0000101101101011";
        wait for clk_period;
        A <= "0001011100001011";
        B <= "0100100001111001";
        C <= "0100011010101111";
        wait for clk_period;
        A <= "1011011100100111";
        B <= "1101000010011100";
        C <= "1100011100010001";
        wait for clk_period;
        A <= "0001001011000001";
        B <= "0000010111110011";
        C <= "0101100111101001";
        wait for clk_period;
        A <= "1111011011110101";
        B <= "0001100111101000";
        C <= "0101001010001001";
        wait for clk_period;
        A <= "1111101111100010";
        B <= "0111100011011100";
        C <= "1000000001000011";
        wait for clk_period;
        A <= "1111011111100100";
        B <= "1011001100110010";
        C <= "1011110011100001";
        wait for clk_period;
        A <= "0000011111111110";
        B <= "0000111001111001";
        C <= "0001001010111100";
        wait for clk_period;
        A <= "0101000011010010";
        B <= "1110001011110100";
        C <= "0101111001011010";
        wait for clk_period;
        A <= "0111110000110001";
        B <= "0111010001011001";
        C <= "1001011111100011";
        wait for clk_period;
        A <= "1110110000000001";
        B <= "0101111100100000";
        C <= "1110000000000001";
        wait for clk_period;
        A <= "1001011000111101";
        B <= "0011010111000110";
        C <= "1010111110000111";
        wait for clk_period;
        A <= "1010101110101100";
        B <= "1110000110011111";
        C <= "1010100010000100";
        wait for clk_period;
        A <= "0000110111111000";
        B <= "0100101101101101";
        C <= "0001110001001101";
        wait for clk_period;
        A <= "1001100011101110";
        B <= "1010110000001001";
        C <= "1001000011000111";
        wait for clk_period;
        A <= "1010010010010001";
        B <= "0111010010011111";
        C <= "1011111000100001";
        wait for clk_period;
        A <= "1000000011111110";
        B <= "0011101011010100";
        C <= "0110100001010101";
        wait for clk_period;
        A <= "0000110100101100";
        B <= "1010011110010111";
        C <= "1000101111011001";
        wait for clk_period;
        A <= "0011011010100010";
        B <= "0110100111000100";
        C <= "0100100000111110";
        wait for clk_period;
        A <= "0101001001111000";
        B <= "1001010101100000";
        C <= "0000010001001001";
        wait for clk_period;
        A <= "1110101010011111";
        B <= "1111010000011101";
        C <= "0011010010111010";
        wait for clk_period;
        A <= "1100001010100101";
        B <= "0111001010100101";
        C <= "1110011010000011";
        wait for clk_period;
        A <= "1000001000111000";
        B <= "0010001101111000";
        C <= "1100101001100110";
        wait for clk_period;
        A <= "0001010001011110";
        B <= "1101011100000000";
        C <= "0101000101111011";
        wait for clk_period;
        A <= "1011010000110110";
        B <= "0101011111100011";
        C <= "1100101110110100";
        wait for clk_period;
        A <= "0011000000001001";
        B <= "0011001111010110";
        C <= "0101110100010110";
        wait for clk_period;
        A <= "0010100010001101";
        B <= "0110111110101011";
        C <= "1110110011111010";
        wait for clk_period;
        A <= "0000001000100101";
        B <= "0100001001110101";
        C <= "0001011000100100";
        wait for clk_period;
        A <= "1100101111001011";
        B <= "1110101101011000";
        C <= "0100011011011010";
        wait for clk_period;
        A <= "0011111001011000";
        B <= "1100100010000000";
        C <= "0100001101111000";
        wait for clk_period;
        A <= "0001110111011011";
        B <= "1101011111101111";
        C <= "1001100011101001";
        wait for clk_period;
        A <= "0000100101101011";
        B <= "1111100100100110";
        C <= "1000101001100011";
        wait for clk_period;
        A <= "0001101101001000";
        B <= "0111010010100100";
        C <= "1110010010000110";
        wait for clk_period;
        A <= "1001110111111011";
        B <= "0111101110111111";
        C <= "0001011011001110";
        wait for clk_period;
        A <= "0000110011011010";
        B <= "1110001101110001";
        C <= "1100111111001100";
        wait for clk_period;
        A <= "0111001011111101";
        B <= "1111100101111111";
        C <= "0111010101100111";
        wait for clk_period;
        A <= "1011001101001000";
        B <= "0101110001010110";
        C <= "1010000111010100";
        wait for clk_period;
        A <= "0111110100100011";
        B <= "0100111101101110";
        C <= "1100101010010010";
        wait for clk_period;
        A <= "0110010000011100";
        B <= "0000100101100110";
        C <= "1001000100110101";
        wait for clk_period;
        A <= "0110001101011101";
        B <= "0101111111101010";
        C <= "1101111000101101";
        wait for clk_period;
        A <= "1101000000101011";
        B <= "1110111110100111";
        C <= "1100000101010011";
        wait for clk_period;
        A <= "1000100001000000";
        B <= "1110000110010000";
        C <= "1111001000110101";
        wait for clk_period;
        A <= "0100111000101100";
        B <= "0011100010000010";
        C <= "0010001010011110";
        wait for clk_period;
        A <= "1000010100001100";
        B <= "0101110011000101";
        C <= "0100011010000000";
        wait for clk_period;
        A <= "1001001010110111";
        B <= "0101100111111110";
        C <= "1011110000001010";
        wait for clk_period;
        A <= "0010001000100100";
        B <= "0110001110011000";
        C <= "0000111101111100";
        wait for clk_period;
        A <= "0010101100011010";
        B <= "1011100001100001";
        C <= "0111111000100010";
        wait for clk_period;
        A <= "1001010101111100";
        B <= "0111110110010111";
        C <= "1000101010001100";
        wait for clk_period;
        A <= "0001100001000111";
        B <= "1000100010110110";
        C <= "1000000011101101";
        wait for clk_period;
        A <= "0011111000000010";
        B <= "0010100001111100";
        C <= "0110010100011101";
        wait for clk_period;
        A <= "1011111111010000";
        B <= "0110000000111011";
        C <= "0000011011001000";
        wait for clk_period;
        A <= "0010101010100111";
        B <= "1000101001010010";
        C <= "1111011100011111";
        wait for clk_period;
        A <= "1110111010000000";
        B <= "0110011111111011";
        C <= "0010011101111000";
        wait for clk_period;
        A <= "0111001100100100";
        B <= "1110000100100010";
        C <= "0000100010010100";
        wait for clk_period;
        A <= "0000000010100110";
        B <= "1001010100011000";
        C <= "1000101011000011";
        wait for clk_period;
        A <= "1011001011111101";
        B <= "1100001010001100";
        C <= "0111101111111000";
        wait for clk_period;
        A <= "1000111110110001";
        B <= "0001111010110011";
        C <= "0010011000111001";
        wait for clk_period;
        A <= "1100001001001001";
        B <= "0011000011001010";
        C <= "1110001001010111";
        wait for clk_period;
        A <= "1111011000010010";
        B <= "1010011010000110";
        C <= "1111000001100111";
        wait for clk_period;
        A <= "1010011010100000";
        B <= "0000010011000011";
        C <= "0000100010101001";
        wait for clk_period;
        A <= "1100110011110011";
        B <= "0000010111100011";
        C <= "1010010100001110";
        wait for clk_period;
        A <= "1010101101110000";
        B <= "1110000001001101";
        C <= "1111011011100011";
        wait for clk_period;
        A <= "0101101111011100";
        B <= "0101010100001101";
        C <= "0011111001101010";
        wait for clk_period;
        A <= "0101011101101100";
        B <= "1100001100101000";
        C <= "0001000000010111";
        wait for clk_period;
        A <= "0001101101111111";
        B <= "1111000011101010";
        C <= "0000010011101001";
        wait for clk_period;
        A <= "1100001101101110";
        B <= "1001010011000011";
        C <= "0110101000010010";
        wait for clk_period;
        A <= "1001111111100011";
        B <= "1001010011111100";
        C <= "0100011011111101";
        wait for clk_period;
        A <= "0110010010100011";
        B <= "0110110011000010";
        C <= "1100000010110111";
        wait for clk_period;
        A <= "0001000110011110";
        B <= "0111111111011101";
        C <= "0101100011111000";
        wait for clk_period;
        A <= "1000111000101101";
        B <= "1011011001011101";
        C <= "1100101011101000";
        wait for clk_period;
        A <= "1000000111111111";
        B <= "1111100100111001";
        C <= "0010111000100101";
        wait for clk_period;
        A <= "0111010111100000";
        B <= "1110010100011100";
        C <= "1001100000011010";
        wait for clk_period;
        A <= "0110100000011001";
        B <= "0111100110001101";
        C <= "1100101000111111";
        wait for clk_period;
        A <= "1011111111100001";
        B <= "1010101011101001";
        C <= "1101111010110101";
        wait for clk_period;
        A <= "0110101101111011";
        B <= "1010111100001101";
        C <= "1000000100001110";
        wait for clk_period;
        A <= "0110011001101101";
        B <= "1111001001011111";
        C <= "1000111100111011";
        wait for clk_period;
        A <= "1110111000010000";
        B <= "1101010001111000";
        C <= "0111101001011010";
        wait for clk_period;
        A <= "1100110011101001";
        B <= "1111110110000001";
        C <= "0100011111111011";
        wait for clk_period;
        A <= "0000000110100111";
        B <= "0100011101011011";
        C <= "0001001010110000";
        wait for clk_period;
        A <= "1100000111101010";
        B <= "0010000100100001";
        C <= "1101110010010011";
        wait for clk_period;
        A <= "0111110011001001";
        B <= "0000101111110010";
        C <= "0100111000100111";
        wait for clk_period;
        A <= "0111001100010011";
        B <= "0001110011111010";
        C <= "0001100010110101";
        wait for clk_period;
        A <= "0001001111011011";
        B <= "0111110000010100";
        C <= "0010011111000000";
        wait for clk_period;
        A <= "1100101101011110";
        B <= "1010101100101100";
        C <= "1111111101110001";
        wait for clk_period;
        A <= "1101101011001001";
        B <= "1100001101100101";
        C <= "1100101011010010";
        wait for clk_period;
        A <= "0011000111100001";
        B <= "0111110100101100";
        C <= "0000011010100010";
        wait for clk_period;
        A <= "1000100010011010";
        B <= "0110010001100111";
        C <= "1101111111101111";
        wait for clk_period;
        A <= "0010000001001110";
        B <= "0111100100111100";
        C <= "1110110111000011";
        wait for clk_period;
        A <= "0011101110010111";
        B <= "1100000010111100";
        C <= "0101001101101101";
        wait for clk_period;
        A <= "0011101111110001";
        B <= "1101101001111001";
        C <= "0000110101001101";
        wait for clk_period;
        A <= "0111000010000000";
        B <= "1110101000010110";
        C <= "0011001011111101";
        wait for clk_period;
        A <= "1011010010000101";
        B <= "0110010010000010";
        C <= "1011010100111000";
        wait for clk_period;
        A <= "1100010011011100";
        B <= "1110100001110000";
        C <= "1010000000100000";
        wait for clk_period;
        A <= "0111111100100001";
        B <= "1110011111111111";
        C <= "0101001001111001";
        wait for clk_period;
        A <= "1110101001000001";
        B <= "0111101010100010";
        C <= "0101011111101100";
        wait for clk_period;
        A <= "1110111000010000";
        B <= "1000101111101000";
        C <= "1110101011110011";
        wait for clk_period;
        A <= "0100011010100011";
        B <= "0000010110111111";
        C <= "1101101110111000";
        wait for clk_period;
        A <= "0010000110110101";
        B <= "1101000010101100";
        C <= "1101101000110111";
        wait for clk_period;
        A <= "1011111010011111";
        B <= "0000010110100011";
        C <= "0110101100010011";
        wait for clk_period;
        A <= "1000110010011111";
        B <= "1111111101001001";
        C <= "1100111101110010";
        wait for clk_period;
        A <= "0100001110011101";
        B <= "1011011001001110";
        C <= "1101000010001001";
        wait for clk_period;
        A <= "0001001110000111";
        B <= "1111101010101000";
        C <= "0101001110000101";
        wait for clk_period;
        A <= "0000101010110001";
        B <= "1000000101001100";
        C <= "1011111100010110";
        wait for clk_period;
        A <= "1101000100011110";
        B <= "0100001111011001";
        C <= "1101001000100001";
        wait for clk_period;
        A <= "1110010100010111";
        B <= "1011000110011100";
        C <= "1000100101000111";
        wait for clk_period;
        A <= "1000101010100010";
        B <= "1011001010111110";
        C <= "1011101101001011";
        wait for clk_period;
        A <= "1011100001000000";
        B <= "1110110100110100";
        C <= "0100110110110100";
        wait for clk_period;
        A <= "0000100011111101";
        B <= "0010011111110000";
        C <= "1001110100011011";
        wait for clk_period;
        A <= "0010100100110000";
        B <= "0111010000011010";
        C <= "1001101001100000";
        wait for clk_period;
        A <= "0101001100011101";
        B <= "1100011111011111";
        C <= "0100011101010111";
        wait for clk_period;
        A <= "1010011101100100";
        B <= "0110101011110101";
        C <= "0100100111001100";
        wait for clk_period;
        A <= "1101011011001101";
        B <= "1000001110101101";
        C <= "1101000000110001";
        wait for clk_period;
        A <= "1101010001001101";
        B <= "0010000010111101";
        C <= "0101010010000000";
        wait for clk_period;
        A <= "1100001100001011";
        B <= "1111011001100000";
        C <= "0101001001100100";
        wait for clk_period;
        A <= "0001000110000001";
        B <= "0101001110101000";
        C <= "1001110000010011";
        wait for clk_period;
        A <= "1000011110011001";
        B <= "0001010000101100";
        C <= "1110011101111011";
        wait for clk_period;
        A <= "0100001100111111";
        B <= "0010110000001001";
        C <= "1101101010000110";
        wait for clk_period;
        A <= "0101000001011100";
        B <= "1010000100001011";
        C <= "0111101010111111";
        wait for clk_period;
        A <= "1010011010011000";
        B <= "1010100001111011";
        C <= "1000011110011101";
        wait for clk_period;
        A <= "1011011101001011";
        B <= "0000000100111001";
        C <= "0110000011001000";
        wait for clk_period;
        A <= "0111000000110100";
        B <= "0111101001111100";
        C <= "0110100001000010";
        wait for clk_period;
        A <= "1110011111001111";
        B <= "1010101011110100";
        C <= "1011100001011101";
        wait for clk_period;
        A <= "1101000000100101";
        B <= "1011100101011110";
        C <= "1100001001010011";
        wait for clk_period;
        A <= "0111001100011110";
        B <= "0011111111011110";
        C <= "1000100000111111";
        wait for clk_period;
        A <= "1010010110000100";
        B <= "1111000110111000";
        C <= "1010100011001001";
        wait for clk_period;
        A <= "1111011110101011";
        B <= "1010010011100111";
        C <= "0111111110011111";
        wait for clk_period;
        A <= "1010111110101100";
        B <= "0100001101011111";
        C <= "0001110100001110";
        wait for clk_period;
        A <= "0100011101110100";
        B <= "0100111101110010";
        C <= "0000000001111111";
        wait for clk_period;
        A <= "1100001011111110";
        B <= "0100101100100100";
        C <= "1010111000001011";
        wait for clk_period;
        A <= "0100011001100111";
        B <= "0010110010111101";
        C <= "1101100000100000";
        wait for clk_period;
        A <= "0111111011101110";
        B <= "0111111011111101";
        C <= "1011110000011110";
        wait for clk_period;
        A <= "0101111101001101";
        B <= "1000111001100000";
        C <= "1001011010100100";
        wait for clk_period;
        A <= "1001010110010100";
        B <= "0110110110000011";
        C <= "0110000001000111";
        wait for clk_period;
        A <= "1011001100110101";
        B <= "1010001010100011";
        C <= "0101110011011000";
        wait for clk_period;
        A <= "0110110111000010";
        B <= "0101000001110011";
        C <= "1100010001011101";
        wait for clk_period;
        A <= "0111101000101110";
        B <= "0101000101100011";
        C <= "0110101110001011";
        wait for clk_period;
        A <= "0001001000101111";
        B <= "0011011000000000";
        C <= "1101010110100111";
        wait for clk_period;
        A <= "0101101001100100";
        B <= "1101010110000110";
        C <= "1110101010011111";
        wait for clk_period;
        A <= "0111001001011011";
        B <= "0100111111001100";
        C <= "1111011101010000";
        wait for clk_period;
        A <= "0101100100010110";
        B <= "1010110100010110";
        C <= "0010111000101101";
        wait for clk_period;
        A <= "1001101000000110";
        B <= "0101100100011001";
        C <= "0100100011100111";
        wait for clk_period;
        A <= "1100110001100111";
        B <= "1000011101001001";
        C <= "1101101001110000";
        wait for clk_period;
        A <= "1111011001111011";
        B <= "0101111010011010";
        C <= "1101101100001111";
        wait for clk_period;
        A <= "1000110100100110";
        B <= "1000001010001111";
        C <= "1100001000001110";
        wait for clk_period;
        A <= "0010110101000001";
        B <= "0110101111100000";
        C <= "1110100110101001";
        wait for clk_period;
        A <= "0011111010001100";
        B <= "1110100111000001";
        C <= "1100010101011100";
        wait for clk_period;
        A <= "0100000011100100";
        B <= "1111010110001110";
        C <= "0001010100101000";
        wait for clk_period;
        A <= "1011100110111010";
        B <= "0011001101110000";
        C <= "1111001000110011";
        wait for clk_period;
        A <= "1001000001101000";
        B <= "1010111001100011";
        C <= "0111001111101100";
        wait for clk_period;
        A <= "0011011111101101";
        B <= "1110010000101011";
        C <= "0100100101010000";
        wait for clk_period;
        A <= "0000111001100110";
        B <= "1010100111110010";
        C <= "0101011110110011";
        wait for clk_period;
        A <= "1001010011000101";
        B <= "1111111010110011";
        C <= "0110010010000001";
        wait for clk_period;
        A <= "1110111101001010";
        B <= "0011101010000101";
        C <= "1001110001000010";
        wait for clk_period;
        A <= "1011011011110011";
        B <= "0000100110000010";
        C <= "1001000101110011";
        wait for clk_period;
        A <= "1000100011110101";
        B <= "0101010001110101";
        C <= "0011110011011111";
        wait for clk_period;
        A <= "0101101000111001";
        B <= "0011101111011010";
        C <= "0010011100110110";
        wait for clk_period;
        A <= "1010001000011001";
        B <= "0011100010100101";
        C <= "0011110101010101";
        wait for clk_period;
        A <= "0011010110111001";
        B <= "0101001110111000";
        C <= "0011010010010110";
        wait for clk_period;
        A <= "0001101000000110";
        B <= "0101101110011010";
        C <= "0011000010100110";
        wait for clk_period;
        A <= "1110100011111101";
        B <= "0100000011011011";
        C <= "0001110110001110";
        wait for clk_period;
        A <= "0111111000000110";
        B <= "0001000000111111";
        C <= "0110101111001100";
        wait for clk_period;
        A <= "1001001111010110";
        B <= "0101001100100011";
        C <= "0000100110111110";
        wait for clk_period;
        A <= "1101001011010111";
        B <= "0000011010100111";
        C <= "0001011000010100";
        wait for clk_period;
        A <= "1010101110001011";
        B <= "1110000010000000";
        C <= "0010101011000101";
        wait for clk_period;
        A <= "1100001001011000";
        B <= "1000100000100111";
        C <= "0011111010000000";
        wait for clk_period;
        A <= "1100101011000111";
        B <= "0100010101011001";
        C <= "0100100100001110";
        wait for clk_period;
        A <= "0010001011010010";
        B <= "1100100101000000";
        C <= "0001000100000110";
        wait for clk_period;
        A <= "0110100110011001";
        B <= "1101110010000110";
        C <= "1011111001100001";
        wait for clk_period;
        A <= "0010101001011010";
        B <= "0011011001101011";
        C <= "0100001011000011";
        wait for clk_period;
        A <= "1101101111001001";
        B <= "0101110001100101";
        C <= "0110111110010000";
        wait for clk_period;
        A <= "1100001010101101";
        B <= "1000001110010101";
        C <= "0111000111011110";
        wait for clk_period;
        A <= "0000001100001110";
        B <= "0010101010100110";
        C <= "0000110001100110";
        wait for clk_period;
        A <= "1101001001010001";
        B <= "0010110010010101";
        C <= "0011110011110110";
        wait for clk_period;
        A <= "0000010100000011";
        B <= "0010001111110010";
        C <= "0110000101110000";
        wait for clk_period;
        A <= "1011111011010011";
        B <= "1000001010110100";
        C <= "1010101001001000";
        wait for clk_period;
        A <= "0100010101110000";
        B <= "0001100111000111";
        C <= "1001001011001001";
        wait for clk_period;
        A <= "1100011011000010";
        B <= "1101000001101111";
        C <= "1110000001011001";
        wait for clk_period;
        A <= "1111011100110101";
        B <= "1000110010001100";
        C <= "0100110011111010";
        wait for clk_period;
        A <= "1110110100001111";
        B <= "0111101010010011";
        C <= "0000111110010011";
        wait for clk_period;
        A <= "1010101110000110";
        B <= "0111001001000011";
        C <= "1111110111010000";
        wait for clk_period;
        A <= "1110111110101011";
        B <= "0100111000010000";
        C <= "0110001101001110";
        wait for clk_period;
        A <= "0001110001011101";
        B <= "1100100001010100";
        C <= "0010010001011010";
        wait for clk_period;
        A <= "0000111011101010";
        B <= "0001111111011000";
        C <= "1000110100111100";
        wait for clk_period;
        A <= "1110001001100101";
        B <= "0101100011101110";
        C <= "0111111000101110";
        wait for clk_period;
        A <= "0110100001001010";
        B <= "1110110011111011";
        C <= "0001011000100011";
        wait for clk_period;
        A <= "0000101001010001";
        B <= "1100101100101011";
        C <= "0110101010110011";
        wait for clk_period;
        A <= "0000001110110100";
        B <= "0100100001010100";
        C <= "0010000100101001";
        wait for clk_period;
        A <= "1011000100010000";
        B <= "0000111000100110";
        C <= "0010001001110001";
        wait for clk_period;
        A <= "1000101101000000";
        B <= "1110001100011101";
        C <= "0001110111010001";
        wait for clk_period;
        A <= "0000100001110011";
        B <= "1001111000010011";
        C <= "1011110110011001";
        wait for clk_period;
        A <= "1110111000001000";
        B <= "1011000001101101";
        C <= "1100000001000010";
        wait for clk_period;
        A <= "1110100010001011";
        B <= "0111101010000011";
        C <= "1010110000111100";
        wait for clk_period;
        A <= "0011111000000000";
        B <= "1111101010010011";
        C <= "0110100100111010";
        wait for clk_period;
        A <= "1111100111001101";
        B <= "1011110000001101";
        C <= "0100010001111011";
        wait for clk_period;
        A <= "1101111111110100";
        B <= "1011101010101101";
        C <= "1011110111000001";
        wait for clk_period;
        A <= "0010101111100011";
        B <= "1111011010001101";
        C <= "0010101110101100";
        wait for clk_period;
        A <= "1101111111000010";
        B <= "0110100110101011";
        C <= "1000001111101100";
        wait for clk_period;
        A <= "1010000111110001";
        B <= "1001110010101110";
        C <= "0101100001101101";
        wait for clk_period;
        A <= "1011100001101100";
        B <= "0010110011000100";
        C <= "1011001001101100";
        wait for clk_period;
        A <= "1010010110010000";
        B <= "1011110100010111";
        C <= "0100101101010010";
        wait for clk_period;
        A <= "1001110111110100";
        B <= "0100101110011111";
        C <= "0100001110000011";
        wait for clk_period;
        A <= "1100111111011101";
        B <= "1001011011111101";
        C <= "0110110100010100";
        wait for clk_period;
        A <= "1001010101100000";
        B <= "0110011001101101";
        C <= "1011100110011110";
        wait for clk_period;
        A <= "0011100101011011";
        B <= "1011110000000110";
        C <= "1101100000110001";
        wait for clk_period;
        A <= "1111011000110100";
        B <= "0001010110100110";
        C <= "0000011001010000";
        wait for clk_period;
        A <= "1010010111011011";
        B <= "1001101011011100";
        C <= "0101001000110100";
        wait for clk_period;
        A <= "0000100100011010";
        B <= "1010100111010100";
        C <= "1000100100001010";
        wait for clk_period;
        A <= "0010001101010101";
        B <= "0101001101111001";
        C <= "0001111000000001";
        wait for clk_period;
        A <= "0011011111000111";
        B <= "1011111101000101";
        C <= "1000011000011011";
        wait for clk_period;
        A <= "0101101101010001";
        B <= "1010001101101111";
        C <= "0111111001100011";
        wait for clk_period;
        A <= "0011001101101101";
        B <= "1111111001100100";
        C <= "1001101001101001";
        wait for clk_period;
        A <= "1110111111011001";
        B <= "0111010011111001";
        C <= "1111011000110100";
        wait for clk_period;
        A <= "1001100001110100";
        B <= "0100001001010001";
        C <= "1100111000101000";
        wait for clk_period;
        A <= "0010010000010010";
        B <= "1001001110111101";
        C <= "0100100010000000";
        wait for clk_period;
        A <= "0000010111001110";
        B <= "0110100000010001";
        C <= "0010011010110010";
        wait for clk_period;
        A <= "0010101011101011";
        B <= "0000100100101001";
        C <= "0011111011111110";
        wait for clk_period;
        A <= "0000010111001110";
        B <= "1110100000101000";
        C <= "0101000011101110";
        wait for clk_period;
        A <= "1111011100100101";
        B <= "0110010000000001";
        C <= "1010000011010000";
        wait for clk_period;
        A <= "0000001101111110";
        B <= "1000001001111010";
        C <= "1001011010101001";
        wait for clk_period;
        A <= "1010110101111111";
        B <= "1001001110000000";
        C <= "1100001110000100";
        wait for clk_period;
        A <= "1001100010101110";
        B <= "0001100100011101";
        C <= "1110001001011011";
        wait for clk_period;
        A <= "1010011110100101";
        B <= "0001001011000010";
        C <= "1101100101011000";
        wait for clk_period;
        A <= "0110101100010010";
        B <= "1101111011010100";
        C <= "1111000101010000";
        wait for clk_period;
        A <= "1000010001011110";
        B <= "1011100000110111";
        C <= "0001100000101100";
        wait for clk_period;
        A <= "1011100111111110";
        B <= "0000010000110101";
        C <= "0111000100010001";
        wait for clk_period;
        A <= "0111011010100110";
        B <= "0101101001100001";
        C <= "1000001011111110";
        wait for clk_period;
        A <= "1011101100000000";
        B <= "0111011111000100";
        C <= "0111000010010010";
        wait for clk_period;
        A <= "1010010111010010";
        B <= "1110000001111001";
        C <= "1101100111010011";
        wait for clk_period;
        A <= "1101101011000100";
        B <= "1100011110110111";
        C <= "0010101001111010";
        wait for clk_period;
        A <= "1001101101010111";
        B <= "1100111100111010";
        C <= "0110100110111111";
        wait for clk_period;
        A <= "1110101100110111";
        B <= "0001011100111110";
        C <= "0011111101100011";
        wait for clk_period;
        A <= "0001101011110011";
        B <= "1101011101001001";
        C <= "0011111000110101";
        wait for clk_period;
        A <= "0110111010100010";
        B <= "0111101100000001";
        C <= "0011010010111100";
        wait for clk_period;
        A <= "0011000111101101";
        B <= "0111000011010100";
        C <= "1101100101110110";
        wait for clk_period;
        A <= "0011100001111001";
        B <= "1111101101010111";
        C <= "0000100001001111";
        wait for clk_period;
        A <= "1100100011111000";
        B <= "0101011001101000";
        C <= "0010100001111110";
        wait for clk_period;
        A <= "0011101110010101";
        B <= "0011011100100100";
        C <= "0111010011111010";
        wait for clk_period;
        A <= "0010110110000000";
        B <= "1001100111010010";
        C <= "1001000000111101";
        wait for clk_period;
        A <= "1110111111000110";
        B <= "1001001100011110";
        C <= "1011000000011010";
        wait for clk_period;
        A <= "0000000000010010";
        B <= "0101011101011001";
        C <= "1111101010110001";
        wait for clk_period;
        A <= "1101010011001111";
        B <= "1000111100011111";
        C <= "1100011000100000";
        wait for clk_period;
        A <= "0011101010000100";
        B <= "1001110110001101";
        C <= "0010000100101110";
        wait for clk_period;
        A <= "1100100010010010";
        B <= "0110000000100011";
        C <= "1011011110010001";
        wait for clk_period;
        A <= "0110001011001101";
        B <= "1111100100000000";
        C <= "0110010110000011";
        wait for clk_period;
        A <= "1001111110111110";
        B <= "0001111010100101";
        C <= "1011011001010000";
        wait for clk_period;
        A <= "0011011101010011";
        B <= "1000110110101111";
        C <= "0110110111001111";
        wait for clk_period;
        A <= "0110101001100001";
        B <= "1111011011111100";
        C <= "1000010100000011";
        wait for clk_period;
        A <= "0001011011111101";
        B <= "0101011101001100";
        C <= "1000000110111111";
        wait for clk_period;
        A <= "1111111101110100";
        B <= "0101101001110000";
        C <= "0101010010100100";
        wait for clk_period;
        A <= "1011000101101111";
        B <= "0110000110001001";
        C <= "0010110011010101";
        wait for clk_period;
        A <= "1100100100001010";
        B <= "1000000100001100";
        C <= "0101011000000000";
        wait for clk_period;
        A <= "1111000111111100";
        B <= "0111001100001001";
        C <= "1100111001001000";
        wait for clk_period;
        A <= "0110000010010001";
        B <= "1011010001001110";
        C <= "0110100110011110";
        wait for clk_period;
        A <= "0101100111111110";
        B <= "0001010111100000";
        C <= "0101010110001010";
        wait for clk_period;
        A <= "0100010111011100";
        B <= "1000111111100001";
        C <= "0011110001100000";
        wait for clk_period;
        A <= "1111010010101001";
        B <= "1111010000000110";
        C <= "1010000001011110";
        wait for clk_period;
        A <= "1110110110100000";
        B <= "1111110001010110";
        C <= "1001011111111110";
        wait for clk_period;
        A <= "0011111101100001";
        B <= "0001010011010001";
        C <= "1011011010010100";
        wait for clk_period;
        A <= "0111001011001101";
        B <= "1011100011101101";
        C <= "1111111011001001";
        wait for clk_period;
        A <= "1101011011100000";
        B <= "1000010011001000";
        C <= "1111011100010101";
        wait for clk_period;
        A <= "0000110111000011";
        B <= "0110111110010101";
        C <= "1101001000111101";
        wait for clk_period;
        A <= "0111110000001011";
        B <= "0000111101001111";
        C <= "1011010100101000";
        wait for clk_period;
        A <= "1010000100100100";
        B <= "0110011101011101";
        C <= "0111111011110110";
        wait for clk_period;
        A <= "1100011001011111";
        B <= "0001000101000111";
        C <= "0001100110011000";
        wait for clk_period;
        A <= "1101111011100001";
        B <= "0110011111000001";
        C <= "0000010100001011";
        wait for clk_period;
        A <= "0111011110010111";
        B <= "0000101110010111";
        C <= "1101011100110010";
        wait for clk_period;
        A <= "0111101111000001";
        B <= "0011100000011110";
        C <= "1001101011010010";
        wait for clk_period;
        A <= "0011111010000001";
        B <= "1100111001011010";
        C <= "0100111001000101";
        wait for clk_period;
        A <= "1000101101001100";
        B <= "0110001100000001";
        C <= "1001000101010011";
        wait for clk_period;
        A <= "0011011000011100";
        B <= "0100001111101110";
        C <= "1011100100010101";
        wait for clk_period;
        A <= "1010100001101001";
        B <= "1101011001000000";
        C <= "1100011001000001";
        wait for clk_period;
        A <= "0101001110101000";
        B <= "0011011100111101";
        C <= "0010011111001111";
        wait for clk_period;
        A <= "0000100101001000";
        B <= "0011010000100111";
        C <= "1100111000110011";
        wait for clk_period;
        A <= "0111001110110000";
        B <= "0101111000101111";
        C <= "1110010110001110";
        wait for clk_period;
        A <= "1100111110000100";
        B <= "0011010010110101";
        C <= "0111110001100110";
        wait for clk_period;
        A <= "0000111000111101";
        B <= "1001011001110011";
        C <= "1001011111110110";
        wait for clk_period;
        A <= "1001001101110111";
        B <= "1101110000011100";
        C <= "1011000011111110";
        wait for clk_period;
        A <= "1101011010110100";
        B <= "0101110000110100";
        C <= "1011011110000110";
        wait for clk_period;
        A <= "0100100001111100";
        B <= "0101001111101101";
        C <= "0110101001011110";
        wait for clk_period;
        A <= "1111100101001001";
        B <= "1000101001010010";
        C <= "0110001010101010";
        wait for clk_period;
        A <= "1110111000111111";
        B <= "1101000001100110";
        C <= "0001100110101010";
        wait for clk_period;
        A <= "1010001100001110";
        B <= "0100000010011100";
        C <= "1001000011001111";
        wait for clk_period;
        A <= "0101001111010011";
        B <= "0011010110000000";
        C <= "0100010111111010";
        wait for clk_period;
        A <= "1001101011000010";
        B <= "0100000001101110";
        C <= "1011011011110100";
        wait for clk_period;
        A <= "1110011011001001";
        B <= "1011100100011000";
        C <= "1011111010011110";
        wait for clk_period;
        A <= "1100111010000001";
        B <= "1101111101111011";
        C <= "1001001010100010";
        wait for clk_period;
        A <= "1011000000010001";
        B <= "1100100111001010";
        C <= "0000000011110011";
        wait for clk_period;
        A <= "0111001110000001";
        B <= "1111001011100001";
        C <= "1001011000100110";
        wait for clk_period;
        A <= "1111010110101101";
        B <= "0111001111101101";
        C <= "0010010111000011";
        wait for clk_period;
        A <= "1111111110110110";
        B <= "0110011111011000";
        C <= "1010100110100001";
        wait for clk_period;
        A <= "0001111111011110";
        B <= "0001100001000000";
        C <= "1111101010110110";
        wait for clk_period;
        A <= "0100010100110000";
        B <= "0001010010001110";
        C <= "1010101110011101";
        wait for clk_period;
        A <= "1000010001001010";
        B <= "1001111010001000";
        C <= "0100100110001111";
        wait for clk_period;
        A <= "0000100001101011";
        B <= "0111001101111011";
        C <= "1010010110110000";
        wait for clk_period;
        A <= "1101111101110000";
        B <= "1011101010101011";
        C <= "1110010101011011";
        wait for clk_period;
        A <= "1101100001011100";
        B <= "0001010110000000";
        C <= "0111011000101011";
        wait for clk_period;
        A <= "0000011101111100";
        B <= "1111100011101111";
        C <= "0110110100100000";
        wait for clk_period;
        A <= "0110100011000110";
        B <= "1110011000000111";
        C <= "0101100000110110";
        wait for clk_period;
        A <= "1111000111111011";
        B <= "0100110000110111";
        C <= "1010101011001011";
        wait for clk_period;
        A <= "0010100101011110";
        B <= "0011010100100101";
        C <= "1011001011001011";
        wait for clk_period;
        A <= "0000111110001011";
        B <= "0110101101100001";
        C <= "1101101101010101";
        wait for clk_period;
        A <= "1000001101001010";
        B <= "1101111100100100";
        C <= "1111110001110001";
        wait for clk_period;
        A <= "0001110111100111";
        B <= "0111100011101011";
        C <= "1001101101000101";
        wait for clk_period;
        A <= "1011011101100000";
        B <= "1011010110100000";
        C <= "1001010000110000";
        wait for clk_period;
        A <= "1000100100100001";
        B <= "1010101101111001";
        C <= "1111010111101001";
        wait for clk_period;
        A <= "1011001111011101";
        B <= "1101000111111101";
        C <= "1010000111000010";
        wait for clk_period;
        A <= "0000111001100110";
        B <= "1111001011111100";
        C <= "0110111001101010";
        wait for clk_period;
        A <= "0001010111110000";
        B <= "0000000011001000";
        C <= "0110000100111110";
        wait for clk_period;
        A <= "1111000101011100";
        B <= "0010010111100110";
        C <= "0000010011111100";
        wait for clk_period;
        A <= "1101000110000100";
        B <= "1100001011010110";
        C <= "0010011110010010";
        wait for clk_period;
        A <= "0101110101010100";
        B <= "1001000101000111";
        C <= "0110010011010100";
        wait for clk_period;
        A <= "0100111010001011";
        B <= "1111111011100100";
        C <= "0100111010001011";
        wait for clk_period;
        A <= "0100000111000010";
        B <= "0100001011101100";
        C <= "0000111011111111";
        wait for clk_period;
        A <= "1010100110000001";
        B <= "1000111101100000";
        C <= "0000001000101110";
        wait for clk_period;
        A <= "1011100000100101";
        B <= "0101100111101111";
        C <= "1000011001111000";
        wait for clk_period;
        A <= "1101110101001111";
        B <= "1010100110110000";
        C <= "0011111100111111";
        wait for clk_period;
        A <= "0001111010000111";
        B <= "0110001001010010";
        C <= "0100000000110011";
        wait for clk_period;
        A <= "1100101000101001";
        B <= "0011000101111010";
        C <= "0001001110100001";
        wait for clk_period;
        A <= "0011101000101101";
        B <= "1111111011110000";
        C <= "0000010110011100";
        wait for clk_period;
        A <= "0001010100111100";
        B <= "1101000000111011";
        C <= "1010001100010010";
        wait for clk_period;
        A <= "1100100101111101";
        B <= "0011111100001100";
        C <= "0000001111111110";
        wait for clk_period;
        A <= "0111111111011010";
        B <= "0011110100101011";
        C <= "1101011101001011";
        wait for clk_period;
        A <= "1101000111010100";
        B <= "1000111000000000";
        C <= "1111011000001101";
        wait for clk_period;
        A <= "1011001111110110";
        B <= "0010010001001011";
        C <= "0011010000011100";
        wait for clk_period;
        A <= "1110111000100010";
        B <= "0000111011111100";
        C <= "1101101100010100";
        wait for clk_period;
        A <= "0101110011111011";
        B <= "0101101011001111";
        C <= "0110111100001010";
        wait for clk_period;
        A <= "1111010101110110";
        B <= "0010111111000001";
        C <= "1110010110100110";
        wait for clk_period;
        A <= "1010010010000001";
        B <= "1100010000010001";
        C <= "0110111001011110";
        wait for clk_period;
        A <= "0100000011101100";
        B <= "1000110111110000";
        C <= "0000100011101110";
        wait for clk_period;
        A <= "1101101001101011";
        B <= "1000010001011101";
        C <= "1100010000101010";
        wait for clk_period;
        A <= "0001110011111011";
        B <= "0001111000000011";
        C <= "0111010011101111";
        wait for clk_period;
        A <= "0000010101111000";
        B <= "1010010000000101";
        C <= "1011111010001111";
        wait for clk_period;
        A <= "0000010000110011";
        B <= "1001101100111010";
        C <= "1100001101011101";
        wait for clk_period;
        A <= "0101011001110011";
        B <= "1000001111011111";
        C <= "0110110111110111";
        wait for clk_period;
        A <= "0011101001110111";
        B <= "0000000110001110";
        C <= "1101101100110100";
        wait for clk_period;
        A <= "0111110000001010";
        B <= "0111100011000000";
        C <= "0111101010111011";
        wait for clk_period;
        A <= "0101111001101101";
        B <= "1110101110000111";
        C <= "1011011100101010";
        wait for clk_period;
        A <= "1101111001101000";
        B <= "0001110110111011";
        C <= "1100111011011100";
        wait for clk_period;
        A <= "1001111000101100";
        B <= "1101000001001000";
        C <= "0001100111001101";
        wait for clk_period;
        A <= "1000001011010100";
        B <= "1110000010000001";
        C <= "1010111110110010";
        wait for clk_period;
        A <= "0100010001110100";
        B <= "0100011001011100";
        C <= "0000101111100001";
        wait for clk_period;
        A <= "0000001110101010";
        B <= "1011110000000010";
        C <= "1110010101000101";
        wait for clk_period;
        A <= "1110110100001000";
        B <= "1110000100001110";
        C <= "0011000100101001";
        wait for clk_period;
        A <= "0100110100001010";
        B <= "0101010011110010";
        C <= "0000010111000001";
        wait for clk_period;
        A <= "1110011010000110";
        B <= "1110111010011110";
        C <= "1000110001001101";
        wait for clk_period;
        A <= "1100010011001100";
        B <= "0010011110001000";
        C <= "0111010111111110";
        wait for clk_period;
        A <= "1011100010101110";
        B <= "1101011010011000";
        C <= "1011011001001010";
        wait for clk_period;
        A <= "1110100001101011";
        B <= "1001011001110110";
        C <= "0101111000111011";
        wait for clk_period;
        A <= "1100101110111100";
        B <= "1010100100111010";
        C <= "1110110110010000";
        wait for clk_period;
        A <= "0001011111111101";
        B <= "1111100101011011";
        C <= "1010010101010011";
        wait for clk_period;
        A <= "0011111111100110";
        B <= "1010111010101110";
        C <= "1000110000001011";
        wait for clk_period;
        A <= "1100001011011110";
        B <= "0111010000110010";
        C <= "0101100110011000";
        wait for clk_period;
        A <= "1011001111110111";
        B <= "1110111010001011";
        C <= "0101111100101100";
        wait for clk_period;
        A <= "0101110011111111";
        B <= "0111001000011101";
        C <= "1110011111011100";
        wait for clk_period;
        A <= "1000001101101001";
        B <= "1110011001111010";
        C <= "1100001000101111";
        wait for clk_period;
        A <= "0001011011001000";
        B <= "0000001101010110";
        C <= "0110010101101111";
        wait for clk_period;
        A <= "0111110001010101";
        B <= "1011111110110010";
        C <= "1001100001101000";
        wait for clk_period;
        A <= "1010011001011000";
        B <= "0010110111100100";
        C <= "1000000011110100";
        wait for clk_period;
        A <= "1011111110000110";
        B <= "1110111000011011";
        C <= "0100110110000000";
        wait for clk_period;
        A <= "1100110011000111";
        B <= "0011001100000111";
        C <= "0001010010000110";
        wait for clk_period;
        A <= "1010000110000100";
        B <= "1011000110100100";
        C <= "1100011100010100";
        wait for clk_period;
        A <= "1001000011011111";
        B <= "0001100100101110";
        C <= "1001101101100110";
        wait for clk_period;
        A <= "1100010101000010";
        B <= "0010001000110110";
        C <= "0001010100101011";
        wait for clk_period;
        A <= "0000110110111111";
        B <= "1100000001000110";
        C <= "1101010001011000";
        wait for clk_period;
        A <= "1000100000000101";
        B <= "1101011010101010";
        C <= "0110011001100011";
        wait for clk_period;
        A <= "1101011101010100";
        B <= "0110010010001111";
        C <= "0010000000110010";
        wait for clk_period;
        A <= "1011101010100000";
        B <= "0101010001111111";
        C <= "0001001011000011";
        wait for clk_period;
        A <= "1011110001100001";
        B <= "0100101111100100";
        C <= "1101000100010100";
        wait for clk_period;
        A <= "0000001010010101";
        B <= "0010100101101101";
        C <= "1100110111100100";
        wait for clk_period;
        A <= "1011100001000011";
        B <= "0110010011101000";
        C <= "0001100000001111";
        wait for clk_period;
        A <= "1011110110100110";
        B <= "1010010000100001";
        C <= "1000010010001111";
        wait for clk_period;
        A <= "1011101000001000";
        B <= "0100111100011100";
        C <= "0001010101100000";
        wait for clk_period;
        A <= "0101101000100101";
        B <= "1000010011011100";
        C <= "0100101110101110";
        wait for clk_period;
        A <= "0000100001010011";
        B <= "1111100110001011";
        C <= "0001100011100011";
        wait for clk_period;
        A <= "0001110000100011";
        B <= "1101100000001100";
        C <= "1101111011011111";
        wait for clk_period;
        A <= "1101110100101111";
        B <= "1000100000001110";
        C <= "1100011011100111";
        wait for clk_period;
        A <= "1110011100111001";
        B <= "1000101100111111";
        C <= "1100010101010011";
        wait for clk_period;
        A <= "1111000000110011";
        B <= "0110001011001100";
        C <= "0010100100110101";
        wait for clk_period;
        A <= "1000111000001101";
        B <= "0011010000011101";
        C <= "0001111001001010";
        wait for clk_period;
        A <= "0010100101011101";
        B <= "0101010001101000";
        C <= "0101011100000111";
        wait for clk_period;
        A <= "0111111010000111";
        B <= "0110000100101001";
        C <= "0101011111001011";
        wait for clk_period;
        A <= "1100110101110101";
        B <= "0100011010110011";
        C <= "1010010001010111";
        wait for clk_period;
        A <= "1100010111101100";
        B <= "1101101111000000";
        C <= "0110010101001001";
        wait for clk_period;
        A <= "1000001011001001";
        B <= "1111000111010111";
        C <= "1110001011110110";
        wait for clk_period;
        A <= "0000011110111110";
        B <= "1101011100000101";
        C <= "1111001101110000";
        wait for clk_period;
        A <= "0111000101001001";
        B <= "0110111110001000";
        C <= "0100000010111010";
        wait for clk_period;
        A <= "0011001111000010";
        B <= "0100010110011000";
        C <= "0111010001000011";
        wait for clk_period;
        A <= "0110110101101101";
        B <= "0110001001111000";
        C <= "0011010110111111";
        wait for clk_period;
        A <= "0111111101001001";
        B <= "0110001111000101";
        C <= "0001101000000000";
        wait for clk_period;
        wait;   
    end process; 
end Behavioral;