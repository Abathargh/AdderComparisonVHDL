library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TB_CSA is
    generic(width: integer := 8);
end TB_CSA;

architecture Behavioral of TB_CSA is

component CarrySaveAdder is
    Port(
        A, B, C: in std_logic_vector(width - 1 downto 0);
        clk: in std_logic;
        Sum: out std_logic_vector(width + 1 downto 0)
    );    
end component;

signal A, B, C: std_logic_vector(width - 1 downto 0);
signal clk: std_logic;
signal Sum: std_logic_vector(width + 1 downto 0);

constant clk_period: time := 2 ns;

begin
    uut: CarrySaveAdder port map(
        A => A,
        B => B,
        C => C,
        clk => clk,
        Sum => Sum
    );
    
    process begin
        clk <= '0';
        wait for clk_period/2;
        clk <= '1';
        wait for clk_period/2;
    end process;

    process begin
        wait for clk_period;
        A <= "10000110";
        B <= "10101001";
        C <= "01010001";
        wait for clk_period;
        A <= "01111010";
        B <= "00111100";
        C <= "01101110";
        wait for clk_period;
        A <= "10010001";
        B <= "10101110";
        C <= "10000101";
        wait for clk_period;
        A <= "00100101";
        B <= "01000101";
        C <= "10111111";
        wait for clk_period;
        A <= "10110000";
        B <= "10111100";
        C <= "10001000";
        wait for clk_period;
        A <= "00111010";
        B <= "01011000";
        C <= "01101101";
        wait for clk_period;
        A <= "10110100";
        B <= "00100001";
        C <= "10110010";
        wait for clk_period;
        A <= "11010110";
        B <= "00101000";
        C <= "01101000";
        wait for clk_period;
        A <= "00000111";
        B <= "11011101";
        C <= "11001100";
        wait for clk_period;
        A <= "11011000";
        B <= "01100100";
        C <= "10110100";
        wait for clk_period;
        A <= "01110100";
        B <= "00111010";
        C <= "11001101";
        wait for clk_period;
        A <= "10111001";
        B <= "10110001";
        C <= "11110110";
        wait for clk_period;
        A <= "10011000";
        B <= "00001100";
        C <= "11100011";
        wait for clk_period;
        A <= "11100101";
        B <= "01110011";
        C <= "10010011";
        wait for clk_period;
        A <= "10001111";
        B <= "00100111";
        C <= "01000100";
        wait for clk_period;
        A <= "10111110";
        B <= "00101011";
        C <= "10100110";
        wait for clk_period;
        A <= "11000011";
        B <= "10110000";
        C <= "01100011";
        wait for clk_period;
        A <= "10000110";
        B <= "10001110";
        C <= "01101100";
        wait for clk_period;
        A <= "01011111";
        B <= "01110110";
        C <= "00110000";
        wait for clk_period;
        A <= "10110110";
        B <= "10001010";
        C <= "01101011";
        wait for clk_period;
        A <= "01111011";
        B <= "00110101";
        C <= "00101001";
        wait for clk_period;
        A <= "10100111";
        B <= "11001111";
        C <= "00000001";
        wait for clk_period;
        A <= "11000100";
        B <= "01001010";
        C <= "00111010";
        wait for clk_period;
        A <= "00001110";
        B <= "10111010";
        C <= "10011111";
        wait for clk_period;
        A <= "11100010";
        B <= "10110000";
        C <= "11010010";
        wait for clk_period;
        A <= "10010100";
        B <= "11110011";
        C <= "01000101";
        wait for clk_period;
        A <= "00011011";
        B <= "10000101";
        C <= "10101011";
        wait for clk_period;
        A <= "11100111";
        B <= "11000110";
        C <= "11100001";
        wait for clk_period;
        A <= "01101000";
        B <= "10011111";
        C <= "11010110";
        wait for clk_period;
        A <= "10111111";
        B <= "00001010";
        C <= "11101111";
        wait for clk_period;
        A <= "10001100";
        B <= "10100111";
        C <= "01001100";
        wait for clk_period;
        A <= "11011011";
        B <= "01011001";
        C <= "00111000";
        wait for clk_period;
        A <= "10101001";
        B <= "11110001";
        C <= "11000110";
        wait for clk_period;
        A <= "11001000";
        B <= "00100111";
        C <= "10011110";
        wait for clk_period;
        A <= "00111100";
        B <= "01100010";
        C <= "01110110";
        wait for clk_period;
        A <= "00100000";
        B <= "01001010";
        C <= "00101100";
        wait for clk_period;
        A <= "11100000";
        B <= "00001101";
        C <= "10000111";
        wait for clk_period;
        A <= "00001011";
        B <= "00010100";
        C <= "01101101";
        wait for clk_period;
        A <= "10011010";
        B <= "11100101";
        C <= "00111010";
        wait for clk_period;
        A <= "10000111";
        B <= "01000000";
        C <= "00000001";
        wait for clk_period;
        A <= "11000001";
        B <= "01011000";
        C <= "10100000";
        wait for clk_period;
        A <= "01001111";
        B <= "01111010";
        C <= "10011000";
        wait for clk_period;
        A <= "10010111";
        B <= "01110101";
        C <= "01110110";
        wait for clk_period;
        A <= "01001010";
        B <= "00101001";
        C <= "11000111";
        wait for clk_period;
        A <= "01110101";
        B <= "01101101";
        C <= "11101010";
        wait for clk_period;
        A <= "11110000";
        B <= "11111101";
        C <= "01010101";
        wait for clk_period;
        A <= "00110001";
        B <= "10101001";
        C <= "01111111";
        wait for clk_period;
        A <= "10100001";
        B <= "01100000";
        C <= "00111101";
        wait for clk_period;
        A <= "01001010";
        B <= "01000010";
        C <= "01100010";
        wait for clk_period;
        A <= "00100111";
        B <= "11100011";
        C <= "11110000";
        wait for clk_period;
        A <= "10101001";
        B <= "11010000";
        C <= "01100101";
        wait for clk_period;
        A <= "00101110";
        B <= "11110101";
        C <= "01010101";
        wait for clk_period;
        A <= "11010001";
        B <= "00000000";
        C <= "01010011";
        wait for clk_period;
        A <= "10011101";
        B <= "10101110";
        C <= "01111001";
        wait for clk_period;
        A <= "00011010";
        B <= "11001011";
        C <= "01000011";
        wait for clk_period;
        A <= "11010100";
        B <= "10111010";
        C <= "00101010";
        wait for clk_period;
        A <= "10000001";
        B <= "01001000";
        C <= "01010110";
        wait for clk_period;
        A <= "01111110";
        B <= "00011011";
        C <= "01101001";
        wait for clk_period;
        A <= "11000110";
        B <= "10010011";
        C <= "11011010";
        wait for clk_period;
        A <= "01100011";
        B <= "10110001";
        C <= "10001110";
        wait for clk_period;
        A <= "11100111";
        B <= "01010000";
        C <= "11001100";
        wait for clk_period;
        A <= "11101100";
        B <= "10100100";
        C <= "11100001";
        wait for clk_period;
        A <= "01101001";
        B <= "11001100";
        C <= "10010011";
        wait for clk_period;
        A <= "10000101";
        B <= "11111001";
        C <= "10111101";
        wait for clk_period;
        A <= "10110110";
        B <= "10111001";
        C <= "11000000";
        wait for clk_period;
        A <= "11110111";
        B <= "01110101";
        C <= "01011000";
        wait for clk_period;
        A <= "01110011";
        B <= "11000000";
        C <= "00001100";
        wait for clk_period;
        A <= "01101001";
        B <= "10101010";
        C <= "01111101";
        wait for clk_period;
        A <= "01110100";
        B <= "11011001";
        C <= "01111010";
        wait for clk_period;
        A <= "00110111";
        B <= "10100000";
        C <= "11101000";
        wait for clk_period;
        A <= "01101100";
        B <= "10001111";
        C <= "11011001";
        wait for clk_period;
        A <= "11011111";
        B <= "11000011";
        C <= "11000001";
        wait for clk_period;
        A <= "01011011";
        B <= "00110100";
        C <= "01110000";
        wait for clk_period;
        A <= "00110101";
        B <= "11010011";
        C <= "10111100";
        wait for clk_period;
        A <= "11010010";
        B <= "10101010";
        C <= "10001010";
        wait for clk_period;
        A <= "11001001";
        B <= "00101100";
        C <= "10111000";
        wait for clk_period;
        A <= "00101000";
        B <= "00000001";
        C <= "11110010";
        wait for clk_period;
        A <= "01101110";
        B <= "10011010";
        C <= "01011100";
        wait for clk_period;
        A <= "11110000";
        B <= "00110000";
        C <= "01010011";
        wait for clk_period;
        A <= "00000001";
        B <= "01011010";
        C <= "10100111";
        wait for clk_period;
        A <= "00011111";
        B <= "01110010";
        C <= "00110110";
        wait for clk_period;
        A <= "00101110";
        B <= "01011101";
        C <= "00100100";
        wait for clk_period;
        A <= "00010011";
        B <= "11010100";
        C <= "00101010";
        wait for clk_period;
        A <= "10110110";
        B <= "11101010";
        C <= "11000010";
        wait for clk_period;
        A <= "11011001";
        B <= "10011110";
        C <= "10101000";
        wait for clk_period;
        A <= "00011101";
        B <= "01101000";
        C <= "10001111";
        wait for clk_period;
        A <= "10111101";
        B <= "11101001";
        C <= "11000110";
        wait for clk_period;
        A <= "10100010";
        B <= "00101010";
        C <= "01010110";
        wait for clk_period;
        A <= "11110110";
        B <= "10001010";
        C <= "00011100";
        wait for clk_period;
        A <= "00000010";
        B <= "00000100";
        C <= "01100010";
        wait for clk_period;
        A <= "11110101";
        B <= "10100100";
        C <= "10101100";
        wait for clk_period;
        A <= "10100000";
        B <= "01011011";
        C <= "01100110";
        wait for clk_period;
        A <= "11000011";
        B <= "11101011";
        C <= "00100111";
        wait for clk_period;
        A <= "11001010";
        B <= "01110011";
        C <= "10010100";
        wait for clk_period;
        A <= "10110000";
        B <= "11110101";
        C <= "00101010";
        wait for clk_period;
        A <= "00011101";
        B <= "00110100";
        C <= "00111101";
        wait for clk_period;
        A <= "10000010";
        B <= "01000011";
        C <= "00000001";
        wait for clk_period;
        A <= "01110100";
        B <= "01011010";
        C <= "10010000";
        wait for clk_period;
        A <= "01100010";
        B <= "00000010";
        C <= "01001011";
        wait for clk_period;
        A <= "10011001";
        B <= "00000000";
        C <= "10100010";
        wait for clk_period;
        A <= "10111111";
        B <= "01101101";
        C <= "00100111";
        wait for clk_period;
        A <= "01000100";
        B <= "11110001";
        C <= "10001000";
        wait for clk_period;
        A <= "01101101";
        B <= "11111001";
        C <= "00101100";
        wait for clk_period;
        A <= "01111110";
        B <= "10001001";
        C <= "11010000";
        wait for clk_period;
        A <= "11010001";
        B <= "11000110";
        C <= "01010110";
        wait for clk_period;
        A <= "00100000";
        B <= "00100110";
        C <= "10111001";
        wait for clk_period;
        A <= "01110001";
        B <= "10011011";
        C <= "01001010";
        wait for clk_period;
        A <= "00010111";
        B <= "10001101";
        C <= "01110000";
        wait for clk_period;
        A <= "00111101";
        B <= "01111000";
        C <= "10000101";
        wait for clk_period;
        A <= "11111011";
        B <= "01110100";
        C <= "00101011";
        wait for clk_period;
        A <= "11101110";
        B <= "00010010";
        C <= "10100101";
        wait for clk_period;
        A <= "11101011";
        B <= "11000110";
        C <= "11100101";
        wait for clk_period;
        A <= "00011101";
        B <= "01100010";
        C <= "10001001";
        wait for clk_period;
        A <= "11110100";
        B <= "10100100";
        C <= "01011101";
        wait for clk_period;
        A <= "00100100";
        B <= "10010110";
        C <= "00011000";
        wait for clk_period;
        A <= "11001011";
        B <= "01010111";
        C <= "01001111";
        wait for clk_period;
        A <= "10000000";
        B <= "11101010";
        C <= "11010011";
        wait for clk_period;
        A <= "00001001";
        B <= "01101111";
        C <= "00011000";
        wait for clk_period;
        A <= "10010101";
        B <= "11001101";
        C <= "11110010";
        wait for clk_period;
        A <= "11010001";
        B <= "11110011";
        C <= "11100010";
        wait for clk_period;
        A <= "11100011";
        B <= "11000100";
        C <= "11100111";
        wait for clk_period;
        A <= "01110001";
        B <= "10101111";
        C <= "10100101";
        wait for clk_period;
        A <= "10001111";
        B <= "11100011";
        C <= "00000110";
        wait for clk_period;
        A <= "00000011";
        B <= "11100101";
        C <= "01011000";
        wait for clk_period;
        A <= "10010001";
        B <= "10100000";
        C <= "01000100";
        wait for clk_period;
        A <= "11110110";
        B <= "11110111";
        C <= "01100000";
        wait for clk_period;
        A <= "11100011";
        B <= "00110001";
        C <= "01100011";
        wait for clk_period;
        A <= "01100011";
        B <= "11110000";
        C <= "10101100";
        wait for clk_period;
        A <= "01001000";
        B <= "00101001";
        C <= "11110001";
        wait for clk_period;
        A <= "00010001";
        B <= "01011101";
        C <= "11110101";
        wait for clk_period;
        A <= "10101111";
        B <= "10000110";
        C <= "00110111";
        wait for clk_period;
        A <= "00110000";
        B <= "01100101";
        C <= "00100000";
        wait for clk_period;
        A <= "00101001";
        B <= "11111001";
        C <= "11010100";
        wait for clk_period;
        A <= "01001101";
        B <= "00010101";
        C <= "11001001";
        wait for clk_period;
        A <= "11001101";
        B <= "11111101";
        C <= "11100111";
        wait for clk_period;
        A <= "00000100";
        B <= "01110100";
        C <= "11011110";
        wait for clk_period;
        A <= "11111011";
        B <= "10100011";
        C <= "11101010";
        wait for clk_period;
        A <= "00101110";
        B <= "11000000";
        C <= "00111001";
        wait for clk_period;
        A <= "01011001";
        B <= "10011100";
        C <= "01000001";
        wait for clk_period;
        A <= "00010111";
        B <= "11010101";
        C <= "11101101";
        wait for clk_period;
        A <= "00000010";
        B <= "10101001";
        C <= "01101010";
        wait for clk_period;
        A <= "01110110";
        B <= "11111111";
        C <= "11000110";
        wait for clk_period;
        A <= "01101111";
        B <= "00000011";
        C <= "10011010";
        wait for clk_period;
        A <= "01110001";
        B <= "11000111";
        C <= "11001000";
        wait for clk_period;
        A <= "10001000";
        B <= "01101100";
        C <= "00111100";
        wait for clk_period;
        A <= "10111110";
        B <= "10100010";
        C <= "10001011";
        wait for clk_period;
        A <= "10111100";
        B <= "10000101";
        C <= "10110010";
        wait for clk_period;
        A <= "00010000";
        B <= "10001000";
        C <= "10111101";
        wait for clk_period;
        A <= "01010010";
        B <= "10111010";
        C <= "00000001";
        wait for clk_period;
        A <= "10111010";
        B <= "10110111";
        C <= "11100011";
        wait for clk_period;
        A <= "01010000";
        B <= "01000101";
        C <= "11000011";
        wait for clk_period;
        A <= "11111101";
        B <= "10111010";
        C <= "10000100";
        wait for clk_period;
        A <= "11100110";
        B <= "01001100";
        C <= "01000000";
        wait for clk_period;
        A <= "10101011";
        B <= "01010101";
        C <= "01001000";
        wait for clk_period;
        A <= "10001000";
        B <= "11001001";
        C <= "11010000";
        wait for clk_period;
        A <= "11000010";
        B <= "01001011";
        C <= "00110100";
        wait for clk_period;
        A <= "01110100";
        B <= "00111110";
        C <= "00001101";
        wait for clk_period;
        A <= "10111010";
        B <= "11011011";
        C <= "01000101";
        wait for clk_period;
        A <= "01010110";
        B <= "00011011";
        C <= "11011100";
        wait for clk_period;
        A <= "10011111";
        B <= "01001010";
        C <= "00000101";
        wait for clk_period;
        A <= "01110111";
        B <= "11010101";
        C <= "01000111";
        wait for clk_period;
        A <= "10100000";
        B <= "10110100";
        C <= "01010011";
        wait for clk_period;
        A <= "01100101";
        B <= "01110011";
        C <= "11100000";
        wait for clk_period;
        A <= "11011001";
        B <= "00011110";
        C <= "00111010";
        wait for clk_period;
        A <= "10000000";
        B <= "00001010";
        C <= "01101011";
        wait for clk_period;
        A <= "00000101";
        B <= "11010000";
        C <= "00100100";
        wait for clk_period;
        A <= "11100100";
        B <= "01000101";
        C <= "01111010";
        wait for clk_period;
        A <= "11010000";
        B <= "11000110";
        C <= "11001100";
        wait for clk_period;
        A <= "00010011";
        B <= "10111011";
        C <= "01110110";
        wait for clk_period;
        A <= "11001111";
        B <= "11010011";
        C <= "00100100";
        wait for clk_period;
        A <= "10100101";
        B <= "01000100";
        C <= "10101110";
        wait for clk_period;
        A <= "11110000";
        B <= "10011000";
        C <= "00001100";
        wait for clk_period;
        A <= "01001110";
        B <= "10010011";
        C <= "11000110";
        wait for clk_period;
        A <= "00011000";
        B <= "11000100";
        C <= "01000100";
        wait for clk_period;
        A <= "10010110";
        B <= "10010011";
        C <= "01000111";
        wait for clk_period;
        A <= "10110001";
        B <= "11000110";
        C <= "01010111";
        wait for clk_period;
        A <= "00101011";
        B <= "10100110";
        C <= "11111010";
        wait for clk_period;
        A <= "01000101";
        B <= "01010110";
        C <= "10100100";
        wait for clk_period;
        A <= "01111101";
        B <= "10011000";
        C <= "01010010";
        wait for clk_period;
        A <= "01110100";
        B <= "11000101";
        C <= "11010101";
        wait for clk_period;
        A <= "11010011";
        B <= "01101001";
        C <= "11001110";
        wait for clk_period;
        A <= "10001000";
        B <= "00010001";
        C <= "10000100";
        wait for clk_period;
        A <= "01100011";
        B <= "00101001";
        C <= "11100110";
        wait for clk_period;
        A <= "11111111";
        B <= "01100010";
        C <= "11101010";
        wait for clk_period;
        A <= "01011000";
        B <= "11010000";
        C <= "10110100";
        wait for clk_period;
        A <= "01100111";
        B <= "10010110";
        C <= "01011010";
        wait for clk_period;
        A <= "00011001";
        B <= "01010010";
        C <= "00100010";
        wait for clk_period;
        A <= "10110011";
        B <= "10010001";
        C <= "11000000";
        wait for clk_period;
        A <= "01000010";
        B <= "10000001";
        C <= "11011001";
        wait for clk_period;
        A <= "10011011";
        B <= "11010111";
        C <= "11001000";
        wait for clk_period;
        A <= "01001110";
        B <= "11110100";
        C <= "00110001";
        wait for clk_period;
        A <= "01010101";
        B <= "10110111";
        C <= "00110111";
        wait for clk_period;
        A <= "00100100";
        B <= "10011010";
        C <= "10101111";
        wait for clk_period;
        A <= "11101100";
        B <= "10110100";
        C <= "11011011";
        wait for clk_period;
        A <= "00011010";
        B <= "01101101";
        C <= "11100101";
        wait for clk_period;
        A <= "10101011";
        B <= "10010111";
        C <= "10001010";
        wait for clk_period;
        A <= "11001110";
        B <= "00101001";
        C <= "00001010";
        wait for clk_period;
        A <= "10101001";
        B <= "00110100";
        C <= "10000001";
        wait for clk_period;
        A <= "00011100";
        B <= "10100000";
        C <= "11110000";
        wait for clk_period;
        A <= "01110011";
        B <= "10110000";
        C <= "01101100";
        wait for clk_period;
        A <= "11100101";
        B <= "00100000";
        C <= "01010100";
        wait for clk_period;
        A <= "10111100";
        B <= "00000111";
        C <= "00011100";
        wait for clk_period;
        A <= "11110001";
        B <= "01100000";
        C <= "01110011";
        wait for clk_period;
        A <= "00100110";
        B <= "11000000";
        C <= "11101011";
        wait for clk_period;
        A <= "10110000";
        B <= "10101001";
        C <= "11101101";
        wait for clk_period;
        A <= "10001100";
        B <= "01111111";
        C <= "00001111";
        wait for clk_period;
        A <= "10000001";
        B <= "10011001";
        C <= "11000000";
        wait for clk_period;
        A <= "01000110";
        B <= "01001010";
        C <= "10001110";
        wait for clk_period;
        A <= "10110100";
        B <= "01011001";
        C <= "10010101";
        wait for clk_period;
        A <= "01100101";
        B <= "11110010";
        C <= "01010101";
        wait for clk_period;
        A <= "01101110";
        B <= "00110001";
        C <= "10000110";
        wait for clk_period;
        A <= "01111101";
        B <= "00010010";
        C <= "00001001";
        wait for clk_period;
        A <= "10101000";
        B <= "11110011";
        C <= "11011110";
        wait for clk_period;
        A <= "11111011";
        B <= "11101100";
        C <= "00000101";
        wait for clk_period;
        A <= "10101100";
        B <= "10111100";
        C <= "10110111";
        wait for clk_period;
        A <= "00110011";
        B <= "00001011";
        C <= "10011001";
        wait for clk_period;
        A <= "10010101";
        B <= "01010011";
        C <= "01010101";
        wait for clk_period;
        A <= "10101000";
        B <= "10001000";
        C <= "01010011";
        wait for clk_period;
        A <= "10101111";
        B <= "11110111";
        C <= "01000101";
        wait for clk_period;
        A <= "01100010";
        B <= "01000101";
        C <= "11011100";
        wait for clk_period;
        A <= "10100011";
        B <= "01011010";
        C <= "10000101";
        wait for clk_period;
        A <= "01001111";
        B <= "00010110";
        C <= "00101110";
        wait for clk_period;
        A <= "01101010";
        B <= "10010000";
        C <= "00111100";
        wait for clk_period;
        A <= "10011011";
        B <= "10111000";
        C <= "10101011";
        wait for clk_period;
        A <= "11001100";
        B <= "11111001";
        C <= "01010100";
        wait for clk_period;
        A <= "11110101";
        B <= "01001110";
        C <= "00101010";
        wait for clk_period;
        A <= "11101111";
        B <= "00101110";
        C <= "10011001";
        wait for clk_period;
        A <= "10010100";
        B <= "11110010";
        C <= "10101101";
        wait for clk_period;
        A <= "10100010";
        B <= "11110000";
        C <= "01010011";
        wait for clk_period;
        A <= "10001000";
        B <= "11000110";
        C <= "11011111";
        wait for clk_period;
        A <= "00111000";
        B <= "00100000";
        C <= "00010011";
        wait for clk_period;
        A <= "00000001";
        B <= "00101110";
        C <= "01001011";
        wait for clk_period;
        A <= "00110011";
        B <= "01110010";
        C <= "11111011";
        wait for clk_period;
        A <= "11001010";
        B <= "11111000";
        C <= "00011110";
        wait for clk_period;
        A <= "10111000";
        B <= "10110011";
        C <= "11110100";
        wait for clk_period;
        A <= "01011100";
        B <= "00000010";
        C <= "11010100";
        wait for clk_period;
        A <= "01100100";
        B <= "00101011";
        C <= "11111000";
        wait for clk_period;
        A <= "00010000";
        B <= "10111110";
        C <= "00010100";
        wait for clk_period;
        A <= "00010011";
        B <= "00110101";
        C <= "01110110";
        wait for clk_period;
        A <= "00100000";
        B <= "10111110";
        C <= "10111000";
        wait for clk_period;
        A <= "01011101";
        B <= "11000010";
        C <= "00101111";
        wait for clk_period;
        A <= "10111001";
        B <= "11011111";
        C <= "11100110";
        wait for clk_period;
        A <= "10001001";
        B <= "01011101";
        C <= "11000010";
        wait for clk_period;
        A <= "01001001";
        B <= "01010001";
        C <= "10001010";
        wait for clk_period;
        A <= "10100000";
        B <= "11000110";
        C <= "10110111";
        wait for clk_period;
        A <= "10110100";
        B <= "11110111";
        C <= "11111000";
        wait for clk_period;
        A <= "11101010";
        B <= "10000101";
        C <= "11110001";
        wait for clk_period;
        A <= "00011100";
        B <= "10010011";
        C <= "10111111";
        wait for clk_period;
        A <= "11000101";
        B <= "10000100";
        C <= "00110100";
        wait for clk_period;
        A <= "10000100";
        B <= "00001011";
        C <= "00010111";
        wait for clk_period;
        A <= "11010010";
        B <= "10011101";
        C <= "00010000";
        wait for clk_period;
        A <= "01101011";
        B <= "11011101";
        C <= "00001001";
        wait for clk_period;
        A <= "00100111";
        B <= "01000100";
        C <= "10100001";
        wait for clk_period;
        A <= "11110111";
        B <= "10100110";
        C <= "00000101";
        wait for clk_period;
        A <= "01111100";
        B <= "11000110";
        C <= "00001010";
        wait for clk_period;
        A <= "01000111";
        B <= "10101110";
        C <= "11110110";
        wait for clk_period;
        A <= "00011001";
        B <= "00110110";
        C <= "01010001";
        wait for clk_period;
        A <= "10010101";
        B <= "10110101";
        C <= "01011000";
        wait for clk_period;
        A <= "00100001";
        B <= "10001100";
        C <= "00010001";
        wait for clk_period;
        A <= "11101011";
        B <= "10101101";
        C <= "11001001";
        wait for clk_period;
        A <= "11010011";
        B <= "11000100";
        C <= "11010100";
        wait for clk_period;
        A <= "10011110";
        B <= "00110101";
        C <= "11110111";
        wait for clk_period;
        A <= "11100100";
        B <= "01000001";
        C <= "11001100";
        wait for clk_period;
        A <= "00000010";
        B <= "00001100";
        C <= "11001010";
        wait for clk_period;
        A <= "10101000";
        B <= "01000110";
        C <= "00100100";
        wait for clk_period;
        A <= "11000000";
        B <= "00011101";
        C <= "10001001";
        wait for clk_period;
        A <= "00100000";
        B <= "10001010";
        C <= "11111110";
        wait for clk_period;
        A <= "10010111";
        B <= "01110010";
        C <= "01111010";
        wait for clk_period;
        A <= "10011010";
        B <= "00010110";
        C <= "00101100";
        wait for clk_period;
        A <= "10011001";
        B <= "00111111";
        C <= "10101000";
        wait for clk_period;
        A <= "01000001";
        B <= "01111110";
        C <= "00101100";
        wait for clk_period;
        A <= "01001101";
        B <= "01001000";
        C <= "11010011";
        wait for clk_period;
        A <= "11011111";
        B <= "00011010";
        C <= "11100110";
        wait for clk_period;
        A <= "11001111";
        B <= "10010111";
        C <= "01110110";
        wait for clk_period;
        A <= "01101111";
        B <= "01101000";
        C <= "11100011";
        wait for clk_period;
        A <= "11000011";
        B <= "10001010";
        C <= "11000000";
        wait for clk_period;
        A <= "01110100";
        B <= "01001100";
        C <= "11011010";
        wait for clk_period;
        A <= "00111111";
        B <= "01100110";
        C <= "11011100";
        wait for clk_period;
        A <= "01100000";
        B <= "01011011";
        C <= "00111110";
        wait for clk_period;
        A <= "01001000";
        B <= "00010001";
        C <= "01110000";
        wait for clk_period;
        A <= "11100100";
        B <= "00110001";
        C <= "10011110";
        wait for clk_period;
        A <= "01011100";
        B <= "11000010";
        C <= "01101001";
        wait for clk_period;
        A <= "11001101";
        B <= "01110000";
        C <= "11010001";
        wait for clk_period;
        A <= "00111101";
        B <= "10101100";
        C <= "10110001";
        wait for clk_period;
        A <= "01000101";
        B <= "11010111";
        C <= "00010111";
        wait for clk_period;
        A <= "00001010";
        B <= "01001000";
        C <= "00101011";
        wait for clk_period;
        A <= "00101100";
        B <= "00100110";
        C <= "10001000";
        wait for clk_period;
        A <= "11011010";
        B <= "01111010";
        C <= "01011110";
        wait for clk_period;
        A <= "00110100";
        B <= "00111101";
        C <= "01101000";
        wait for clk_period;
        A <= "01110000";
        B <= "01001111";
        C <= "11000001";
        wait for clk_period;
        A <= "00101011";
        B <= "10101100";
        C <= "10110010";
        wait for clk_period;
        A <= "01010001";
        B <= "00001010";
        C <= "01100010";
        wait for clk_period;
        A <= "10110101";
        B <= "11000011";
        C <= "10101011";
        wait for clk_period;
        A <= "01111101";
        B <= "00000001";
        C <= "10011001";
        wait for clk_period;
        A <= "01000111";
        B <= "01001010";
        C <= "11101111";
        wait for clk_period;
        A <= "11011001";
        B <= "00001010";
        C <= "10100111";
        wait for clk_period;
        A <= "10111001";
        B <= "00001010";
        C <= "10110110";
        wait for clk_period;
        A <= "11101001";
        B <= "00011110";
        C <= "00101110";
        wait for clk_period;
        A <= "10000000";
        B <= "10100111";
        C <= "10010111";
        wait for clk_period;
        A <= "00011011";
        B <= "01010010";
        C <= "00011100";
        wait for clk_period;
        A <= "01111100";
        B <= "11101010";
        C <= "00100111";
        wait for clk_period;
        A <= "10001101";
        B <= "11110110";
        C <= "11101000";
        wait for clk_period;
        A <= "10101001";
        B <= "00010011";
        C <= "01110010";
        wait for clk_period;
        A <= "01011111";
        B <= "10101101";
        C <= "00010000";
        wait for clk_period;
        A <= "00010010";
        B <= "10101101";
        C <= "11010001";
        wait for clk_period;
        A <= "00111110";
        B <= "00101111";
        C <= "01111110";
        wait for clk_period;
        A <= "10100011";
        B <= "00010100";
        C <= "00000100";
        wait for clk_period;
        A <= "10111111";
        B <= "10000111";
        C <= "10001010";
        wait for clk_period;
        A <= "00111111";
        B <= "00100010";
        C <= "01110111";
        wait for clk_period;
        A <= "11001101";
        B <= "01001001";
        C <= "11011111";
        wait for clk_period;
        A <= "11111100";
        B <= "00011001";
        C <= "01011101";
        wait for clk_period;
        A <= "00011101";
        B <= "11010100";
        C <= "11101111";
        wait for clk_period;
        A <= "00111001";
        B <= "00110001";
        C <= "00110010";
        wait for clk_period;
        A <= "00000011";
        B <= "11000011";
        C <= "10100110";
        wait for clk_period;
        A <= "11000011";
        B <= "11111011";
        C <= "11110100";
        wait for clk_period;
        A <= "10111011";
        B <= "10011010";
        C <= "01001010";
        wait for clk_period;
        A <= "00000101";
        B <= "10100111";
        C <= "00011010";
        wait for clk_period;
        A <= "01110011";
        B <= "10001010";
        C <= "01011000";
        wait for clk_period;
        A <= "00011100";
        B <= "00101001";
        C <= "01111011";
        wait for clk_period;
        A <= "10100100";
        B <= "01110101";
        C <= "01010100";
        wait for clk_period;
        A <= "11111101";
        B <= "01011000";
        C <= "11011010";
        wait for clk_period;
        A <= "10001001";
        B <= "01010100";
        C <= "11111111";
        wait for clk_period;
        A <= "00111111";
        B <= "00111111";
        C <= "11100010";
        wait for clk_period;
        A <= "11101011";
        B <= "01111110";
        C <= "11111010";
        wait for clk_period;
        A <= "00001001";
        B <= "11000010";
        C <= "11100001";
        wait for clk_period;
        A <= "11000101";
        B <= "00100101";
        C <= "11011001";
        wait for clk_period;
        A <= "01100101";
        B <= "01000010";
        C <= "11010111";
        wait for clk_period;
        A <= "11011111";
        B <= "10101001";
        C <= "01000101";
        wait for clk_period;
        A <= "11010011";
        B <= "10010011";
        C <= "00010010";
        wait for clk_period;
        A <= "01101000";
        B <= "11110110";
        C <= "10010001";
        wait for clk_period;
        A <= "11001001";
        B <= "10010100";
        C <= "01111000";
        wait for clk_period;
        A <= "01001001";
        B <= "11001101";
        C <= "10110001";
        wait for clk_period;
        A <= "11011111";
        B <= "00100000";
        C <= "10011001";
        wait for clk_period;
        A <= "00010011";
        B <= "11111110";
        C <= "01011000";
        wait for clk_period;
        A <= "00100101";
        B <= "01110000";
        C <= "01010111";
        wait for clk_period;
        A <= "00111111";
        B <= "01011101";
        C <= "00010000";
        wait for clk_period;
        A <= "11011000";
        B <= "00001010";
        C <= "00010101";
        wait for clk_period;
        A <= "10011100";
        B <= "01000011";
        C <= "00000101";
        wait for clk_period;
        A <= "10001111";
        B <= "10110000";
        C <= "00010111";
        wait for clk_period;
        A <= "01001110";
        B <= "10110000";
        C <= "01000011";
        wait for clk_period;
        A <= "11001010";
        B <= "01000011";
        C <= "10111100";
        wait for clk_period;
        A <= "10000000";
        B <= "10110010";
        C <= "10110010";
        wait for clk_period;
        A <= "01111001";
        B <= "01101011";
        C <= "01000100";
        wait for clk_period;
        A <= "01010011";
        B <= "10001111";
        C <= "00110110";
        wait for clk_period;
        A <= "10011010";
        B <= "00101010";
        C <= "01001101";
        wait for clk_period;
        A <= "00001110";
        B <= "11110000";
        C <= "01010000";
        wait for clk_period;
        A <= "00100111";
        B <= "11000101";
        C <= "11001101";
        wait for clk_period;
        A <= "01110001";
        B <= "01111110";
        C <= "01000010";
        wait for clk_period;
        A <= "01000100";
        B <= "00110010";
        C <= "11111101";
        wait for clk_period;
        A <= "00010110";
        B <= "10111111";
        C <= "00110111";
        wait for clk_period;
        A <= "00110101";
        B <= "11110010";
        C <= "01111011";
        wait for clk_period;
        A <= "00100010";
        B <= "11011110";
        C <= "11101000";
        wait for clk_period;
        A <= "11000001";
        B <= "11010011";
        C <= "01100000";
        wait for clk_period;
        A <= "10110010";
        B <= "01011111";
        C <= "11000101";
        wait for clk_period;
        A <= "00000011";
        B <= "10111110";
        C <= "00010001";
        wait for clk_period;
        A <= "00110000";
        B <= "11111110";
        C <= "11010100";
        wait for clk_period;
        A <= "10011010";
        B <= "00000100";
        C <= "10111111";
        wait for clk_period;
        A <= "11101101";
        B <= "11010011";
        C <= "01010001";
        wait for clk_period;
        A <= "10110100";
        B <= "11111111";
        C <= "10110000";
        wait for clk_period;
        A <= "11100001";
        B <= "11111000";
        C <= "01110000";
        wait for clk_period;
        A <= "10000111";
        B <= "11100110";
        C <= "00010000";
        wait for clk_period;
        A <= "11110110";
        B <= "00011111";
        C <= "11101001";
        wait for clk_period;
        A <= "11101011";
        B <= "10010110";
        C <= "00101111";
        wait for clk_period;
        A <= "10001000";
        B <= "00010111";
        C <= "11111111";
        wait for clk_period;
        A <= "11010100";
        B <= "11010110";
        C <= "00111111";
        wait for clk_period;
        A <= "10011010";
        B <= "01001110";
        C <= "10001100";
        wait for clk_period;
        A <= "10001000";
        B <= "10011101";
        C <= "01001001";
        wait for clk_period;
        A <= "00011010";
        B <= "01001100";
        C <= "10000101";
        wait for clk_period;
        A <= "10011011";
        B <= "10101100";
        C <= "11111100";
        wait for clk_period;
        A <= "11101001";
        B <= "01001110";
        C <= "01100000";
        wait for clk_period;
        A <= "01111011";
        B <= "10100110";
        C <= "10101100";
        wait for clk_period;
        A <= "00000111";
        B <= "11001010";
        C <= "10111011";
        wait for clk_period;
        A <= "00000000";
        B <= "01011111";
        C <= "10100001";
        wait for clk_period;
        A <= "10010011";
        B <= "00000111";
        C <= "01001100";
        wait for clk_period;
        A <= "00110010";
        B <= "10000110";
        C <= "11010100";
        wait for clk_period;
        A <= "10000100";
        B <= "11101000";
        C <= "01101011";
        wait for clk_period;
        A <= "10001011";
        B <= "01101100";
        C <= "01111101";
        wait for clk_period;
        A <= "00010010";
        B <= "11011010";
        C <= "01110101";
        wait for clk_period;
        A <= "11111100";
        B <= "11010100";
        C <= "11010111";
        wait for clk_period;
        A <= "00100101";
        B <= "00101000";
        C <= "01001001";
        wait for clk_period;
        A <= "00101000";
        B <= "11101111";
        C <= "01000110";
        wait for clk_period;
        A <= "00001000";
        B <= "01011011";
        C <= "01011010";
        wait for clk_period;
        A <= "10001110";
        B <= "00110011";
        C <= "01111100";
        wait for clk_period;
        A <= "11010000";
        B <= "00101010";
        C <= "10000010";
        wait for clk_period;
        A <= "10100000";
        B <= "01010101";
        C <= "01110001";
        wait for clk_period;
        A <= "01110001";
        B <= "00101010";
        C <= "01000101";
        wait for clk_period;
        A <= "01110101";
        B <= "01100110";
        C <= "11110110";
        wait for clk_period;
        A <= "11011100";
        B <= "01101011";
        C <= "00010101";
        wait for clk_period;
        A <= "10101111";
        B <= "00110101";
        C <= "10101010";
        wait for clk_period;
        A <= "01101100";
        B <= "10111000";
        C <= "11000101";
        wait for clk_period;
        A <= "00010000";
        B <= "00111110";
        C <= "11000010";
        wait for clk_period;
        A <= "01100000";
        B <= "10110100";
        C <= "00001010";
        wait for clk_period;
        A <= "00001111";
        B <= "00001101";
        C <= "01100001";
        wait for clk_period;
        A <= "10010111";
        B <= "11110101";
        C <= "01110110";
        wait for clk_period;
        A <= "00011100";
        B <= "01100101";
        C <= "00010011";
        wait for clk_period;
        A <= "01000110";
        B <= "00100100";
        C <= "01101001";
        wait for clk_period;
        A <= "00000111";
        B <= "01001001";
        C <= "11110100";
        wait for clk_period;
        A <= "10111111";
        B <= "10011011";
        C <= "11111111";
        wait for clk_period;
        A <= "01010101";
        B <= "00100000";
        C <= "10010010";
        wait for clk_period;
        A <= "01011011";
        B <= "11010011";
        C <= "10000111";
        wait for clk_period;
        A <= "10001101";
        B <= "10101110";
        C <= "01100110";
        wait for clk_period;
        A <= "11000101";
        B <= "01010010";
        C <= "01110111";
        wait for clk_period;
        A <= "11101010";
        B <= "00011011";
        C <= "00010000";
        wait for clk_period;
        A <= "00011010";
        B <= "00100101";
        C <= "11110110";
        wait for clk_period;
        A <= "10101011";
        B <= "00001101";
        C <= "11010001";
        wait for clk_period;
        A <= "01100011";
        B <= "01100110";
        C <= "01111111";
        wait for clk_period;
        A <= "01111010";
        B <= "11101010";
        C <= "01010010";
        wait for clk_period;
        A <= "00101100";
        B <= "01101000";
        C <= "11111010";
        wait for clk_period;
        A <= "10001000";
        B <= "11110011";
        C <= "10000101";
        wait for clk_period;
        A <= "01110111";
        B <= "01110111";
        C <= "00010100";
        wait for clk_period;
        A <= "01000100";
        B <= "00101011";
        C <= "11010110";
        wait for clk_period;
        A <= "01011000";
        B <= "01000110";
        C <= "00101111";
        wait for clk_period;
        A <= "11010100";
        B <= "10010111";
        C <= "00111010";
        wait for clk_period;
        A <= "01111001";
        B <= "00010110";
        C <= "11111010";
        wait for clk_period;
        A <= "00010000";
        B <= "10001110";
        C <= "00010000";
        wait for clk_period;
        A <= "11010111";
        B <= "01000010";
        C <= "00100101";
        wait for clk_period;
        A <= "00010000";
        B <= "10010010";
        C <= "00101111";
        wait for clk_period;
        A <= "11111001";
        B <= "11010111";
        C <= "10001100";
        wait for clk_period;
        A <= "01111001";
        B <= "10001000";
        C <= "00001010";
        wait for clk_period;
        A <= "01000111";
        B <= "00011011";
        C <= "01100011";
        wait for clk_period;
        A <= "11011001";
        B <= "01110001";
        C <= "00001101";
        wait for clk_period;
        A <= "01110001";
        B <= "11101110";
        C <= "10100000";
        wait for clk_period;
        A <= "10001011";
        B <= "00100100";
        C <= "10001000";
        wait for clk_period;
        A <= "10100011";
        B <= "10011101";
        C <= "00100011";
        wait for clk_period;
        A <= "00100010";
        B <= "11000100";
        C <= "01000001";
        wait for clk_period;
        A <= "10100001";
        B <= "01111010";
        C <= "00101000";
        wait for clk_period;
        A <= "01101011";
        B <= "01100000";
        C <= "01111010";
        wait for clk_period;
        A <= "01010100";
        B <= "11000110";
        C <= "00000100";
        wait for clk_period;
        A <= "00101110";
        B <= "00011001";
        C <= "01010001";
        wait for clk_period;
        A <= "00111011";
        B <= "11100100";
        C <= "10010010";
        wait for clk_period;
        A <= "10001011";
        B <= "01101101";
        C <= "11011100";
        wait for clk_period;
        A <= "01000100";
        B <= "00000101";
        C <= "00111010";
        wait for clk_period;
        A <= "01010110";
        B <= "11101110";
        C <= "01110101";
        wait for clk_period;
        A <= "10010000";
        B <= "10110101";
        C <= "01101111";
        wait for clk_period;
        A <= "00011011";
        B <= "01010110";
        C <= "01100100";
        wait for clk_period;
        A <= "10000000";
        B <= "00111001";
        C <= "01100111";
        wait for clk_period;
        A <= "00110010";
        B <= "11000111";
        C <= "00110110";
        wait for clk_period;
        A <= "10100101";
        B <= "10001011";
        C <= "10110000";
        wait for clk_period;
        A <= "01101111";
        B <= "11010111";
        C <= "00110011";
        wait for clk_period;
        A <= "01010001";
        B <= "00001101";
        C <= "10010110";
        wait for clk_period;
        A <= "11111010";
        B <= "11000011";
        C <= "01111011";
        wait for clk_period;
        A <= "01010011";
        B <= "00101101";
        C <= "10011100";
        wait for clk_period;
        A <= "00111111";
        B <= "11111011";
        C <= "00100000";
        wait for clk_period;
        A <= "11010101";
        B <= "01000000";
        C <= "01001000";
        wait for clk_period;
        A <= "00101110";
        B <= "11111001";
        C <= "10111110";
        wait for clk_period;
        A <= "11001111";
        B <= "00110011";
        C <= "00110110";
        wait for clk_period;
        A <= "00010111";
        B <= "11100110";
        C <= "10110011";
        wait for clk_period;
        A <= "11110110";
        B <= "01110011";
        C <= "11100010";
        wait for clk_period;
        A <= "01111100";
        B <= "00100101";
        C <= "01110010";
        wait for clk_period;
        A <= "11101000";
        B <= "01011011";
        C <= "01000000";
        wait for clk_period;
        A <= "00010001";
        B <= "00111111";
        C <= "00011000";
        wait for clk_period;
        A <= "11010000";
        B <= "11010010";
        C <= "11110100";
        wait for clk_period;
        A <= "01010001";
        B <= "00010101";
        C <= "10101100";
        wait for clk_period;
        A <= "01101011";
        B <= "10011001";
        C <= "00010110";
        wait for clk_period;
        A <= "01111111";
        B <= "11000111";
        C <= "00110000";
        wait for clk_period;
        A <= "00111001";
        B <= "01011000";
        C <= "11110011";
        wait for clk_period;
        A <= "10000100";
        B <= "00011110";
        C <= "00110110";
        wait for clk_period;
        A <= "00011111";
        B <= "10100100";
        C <= "11110000";
        wait for clk_period;
        A <= "10000011";
        B <= "11010111";
        C <= "01010111";
        wait for clk_period;
        A <= "00011101";
        B <= "10101011";
        C <= "11010111";
        wait for clk_period;
        A <= "01111100";
        B <= "00000001";
        C <= "11001111";
        wait for clk_period;
        A <= "01100011";
        B <= "01011110";
        C <= "11001100";
        wait for clk_period;
        A <= "11111011";
        B <= "10111011";
        C <= "01101001";
        wait for clk_period;
        A <= "10010010";
        B <= "10010011";
        C <= "10011101";
        wait for clk_period;
        A <= "01001011";
        B <= "00101001";
        C <= "10001101";
        wait for clk_period;
        A <= "01110101";
        B <= "01010011";
        C <= "11100101";
        wait for clk_period;
        A <= "10011111";
        B <= "10010110";
        C <= "00011001";
        wait for clk_period;
        A <= "01011110";
        B <= "10011101";
        C <= "00110111";
        wait for clk_period;
        A <= "10001100";
        B <= "10100000";
        C <= "01001011";
        wait for clk_period;
        A <= "10101010";
        B <= "00101101";
        C <= "11000000";
        wait for clk_period;
        A <= "01000010";
        B <= "10010100";
        C <= "01000000";
        wait for clk_period;
        A <= "01110011";
        B <= "11000101";
        C <= "10100111";
        wait for clk_period;
        A <= "11010010";
        B <= "11100100";
        C <= "10011001";
        wait for clk_period;
        A <= "10011000";
        B <= "11101101";
        C <= "10010101";
        wait for clk_period;
        A <= "00110011";
        B <= "00001111";
        C <= "01100010";
        wait for clk_period;
        A <= "11100010";
        B <= "10101110";
        C <= "10000100";
        wait for clk_period;
        A <= "11110110";
        B <= "00001111";
        C <= "10011011";
        wait for clk_period;
        A <= "00100110";
        B <= "01100010";
        C <= "00111010";
        wait for clk_period;
        A <= "01001101";
        B <= "01010000";
        C <= "01111000";
        wait for clk_period;
        A <= "01101101";
        B <= "10001110";
        C <= "11111000";
        wait for clk_period;
        A <= "11111101";
        B <= "01110011";
        C <= "01010110";
        wait for clk_period;
        A <= "11101010";
        B <= "11101000";
        C <= "10011101";
        wait for clk_period;
        A <= "01011011";
        B <= "01010010";
        C <= "00000111";
        wait for clk_period;
        A <= "01100100";
        B <= "11011000";
        C <= "01001011";
        wait for clk_period;
        A <= "00100110";
        B <= "11011100";
        C <= "10011100";
        wait for clk_period;
        A <= "00010101";
        B <= "00011110";
        C <= "10010100";
        wait for clk_period;
        A <= "11010101";
        B <= "00010010";
        C <= "01011010";
        wait for clk_period;
        A <= "11100111";
        B <= "00001110";
        C <= "00111101";
        wait for clk_period;
        A <= "01110011";
        B <= "00010110";
        C <= "00010000";
        wait for clk_period;
        A <= "00011010";
        B <= "10000110";
        C <= "10110001";
        wait for clk_period;
        A <= "11000011";
        B <= "00001000";
        C <= "01001011";
        wait for clk_period;
        A <= "01011001";
        B <= "11000111";
        C <= "00111111";
        wait for clk_period;
        A <= "00010000";
        B <= "01011011";
        C <= "00001000";
        wait for clk_period;
        A <= "00110101";
        B <= "11011000";
        C <= "11011110";
        wait for clk_period;
        A <= "11010101";
        B <= "00010000";
        C <= "11111001";
        wait for clk_period;
        A <= "10100011";
        B <= "01000010";
        C <= "01111011";
        wait for clk_period;
        A <= "00000101";
        B <= "10101100";
        C <= "10111011";
        wait for clk_period;
        A <= "00111101";
        B <= "11101011";
        C <= "01110110";
        wait for clk_period;
        A <= "11001000";
        B <= "00100111";
        C <= "00100010";
        wait for clk_period;
        A <= "10100001";
        B <= "11111100";
        C <= "00010011";
        wait for clk_period;
        A <= "01010001";
        B <= "01110110";
        C <= "11011011";
        wait for clk_period;
        A <= "01010100";
        B <= "10100110";
        C <= "00100010";
        wait for clk_period;
        A <= "11101100";
        B <= "01001011";
        C <= "01110010";
        wait for clk_period;
        A <= "01100110";
        B <= "01001111";
        C <= "11110001";
        wait for clk_period;
        A <= "10111010";
        B <= "10011100";
        C <= "10101110";
        wait for clk_period;
        A <= "01000111";
        B <= "11100001";
        C <= "00110010";
        wait for clk_period;
        A <= "01100011";
        B <= "11101010";
        C <= "10100000";
        wait for clk_period;
        A <= "00100001";
        B <= "00100010";
        C <= "01110000";
        wait for clk_period;
        A <= "01010011";
        B <= "00000100";
        C <= "01100110";
        wait for clk_period;
        A <= "00011110";
        B <= "11110111";
        C <= "01110111";
        wait for clk_period;
        A <= "10101101";
        B <= "00110011";
        C <= "01011000";
        wait for clk_period;
        A <= "10110010";
        B <= "11101100";
        C <= "11000110";
        wait for clk_period;
        A <= "10010100";
        B <= "11111101";
        C <= "10000101";
        wait for clk_period;
        A <= "10011011";
        B <= "01111110";
        C <= "00110101";
        wait for clk_period;
        A <= "01001110";
        B <= "00011000";
        C <= "11010100";
        wait for clk_period;
        A <= "00011111";
        B <= "10010000";
        C <= "01011001";
        wait for clk_period;
        A <= "10010011";
        B <= "01110110";
        C <= "10101001";
        wait for clk_period;
        A <= "11111000";
        B <= "01110101";
        C <= "10100000";
        wait for clk_period;
        A <= "01000000";
        B <= "00011111";
        C <= "00111101";
        wait for clk_period;
        A <= "11000010";
        B <= "11011101";
        C <= "00001010";
        wait for clk_period;
        A <= "10110110";
        B <= "10110000";
        C <= "11001101";
        wait for clk_period;
        A <= "10010000";
        B <= "00110010";
        C <= "11010000";
        wait for clk_period;
        A <= "00110001";
        B <= "01101001";
        C <= "11011010";
        wait for clk_period;
        A <= "00110011";
        B <= "01010100";
        C <= "01100110";
        wait for clk_period;
        A <= "00000001";
        B <= "00001001";
        C <= "11110010";
        wait for clk_period;
        A <= "11001000";
        B <= "00101111";
        C <= "11000001";
        wait for clk_period;
        A <= "11100010";
        B <= "01110111";
        C <= "00000011";
        wait for clk_period;
        A <= "10011110";
        B <= "10011100";
        C <= "00010111";
        wait for clk_period;
        A <= "00110000";
        B <= "11010010";
        C <= "10111000";
        wait for clk_period;
        A <= "11100010";
        B <= "00101011";
        C <= "11110110";
        wait for clk_period;
        A <= "01011011";
        B <= "01010001";
        C <= "00110011";
        wait for clk_period;
        A <= "01011000";
        B <= "11110110";
        C <= "11010101";
        wait for clk_period;
        A <= "01110011";
        B <= "01000111";
        C <= "00011010";
        wait for clk_period;
        A <= "00000100";
        B <= "11111000";
        C <= "11110100";
        wait for clk_period;
        A <= "11011110";
        B <= "11000011";
        C <= "10011101";
        wait for clk_period;
        A <= "10011011";
        B <= "10010001";
        C <= "11100110";
        wait for clk_period;
        A <= "00010010";
        B <= "11100000";
        C <= "10000111";
        wait for clk_period;
        A <= "01111001";
        B <= "00111110";
        C <= "01010110";
        wait for clk_period;
        A <= "01011001";
        B <= "01001011";
        C <= "10101110";
        wait for clk_period;
        A <= "10101011";
        B <= "10001100";
        C <= "10110101";
        wait for clk_period;
        A <= "10000111";
        B <= "01001111";
        C <= "11000011";
        wait for clk_period;
        A <= "00011011";
        B <= "10101110";
        C <= "01000010";
        wait for clk_period;
        A <= "10001100";
        B <= "10100000";
        C <= "11110110";
        wait for clk_period;
        A <= "10111110";
        B <= "01000010";
        C <= "01100101";
        wait for clk_period;
        A <= "00001100";
        B <= "00010010";
        C <= "10011010";
        wait for clk_period;
        A <= "01110001";
        B <= "10000000";
        C <= "10010000";
        wait for clk_period;
        A <= "00000000";
        B <= "01100000";
        C <= "00011000";
        wait for clk_period;
        A <= "10101011";
        B <= "10100110";
        C <= "10010011";
        wait for clk_period;
        A <= "00001011";
        B <= "11011000";
        C <= "00101001";
        wait for clk_period;
        A <= "01000000";
        B <= "10010011";
        C <= "11001100";
        wait for clk_period;
        A <= "00010111";
        B <= "01101011";
        C <= "00100001";
        wait for clk_period;
        A <= "01011110";
        B <= "10011111";
        C <= "10000101";
        wait for clk_period;
        A <= "11000010";
        B <= "10001100";
        C <= "11110001";
        wait for clk_period;
        A <= "11000010";
        B <= "10101010";
        C <= "00000010";
        wait for clk_period;
        A <= "11111111";
        B <= "11101101";
        C <= "11010011";
        wait for clk_period;
        A <= "11001000";
        B <= "01001100";
        C <= "00010010";
        wait for clk_period;
        A <= "11010001";
        B <= "10111001";
        C <= "11001101";
        wait for clk_period;
        A <= "11110001";
        B <= "00101001";
        C <= "01010011";
        wait for clk_period;
        A <= "00011010";
        B <= "00000111";
        C <= "00101010";
        wait for clk_period;
        A <= "10101100";
        B <= "00000010";
        C <= "01001000";
        wait for clk_period;
        A <= "11110100";
        B <= "11000111";
        C <= "10001111";
        wait for clk_period;
        A <= "10010000";
        B <= "00110100";
        C <= "10010001";
        wait for clk_period;
        A <= "10100101";
        B <= "11010011";
        C <= "00001101";
        wait for clk_period;
        A <= "11111101";
        B <= "10010010";
        C <= "11111011";
        wait for clk_period;
        A <= "00001010";
        B <= "01001010";
        C <= "01111000";
        wait for clk_period;
        A <= "10110000";
        B <= "00001100";
        C <= "11110101";
        wait for clk_period;
        A <= "00001111";
        B <= "10010011";
        C <= "10100100";
        wait for clk_period;
        A <= "10010000";
        B <= "10010110";
        C <= "11101110";
        wait for clk_period;
        A <= "10100000";
        B <= "01001101";
        C <= "01101100";
        wait for clk_period;
        A <= "00111110";
        B <= "11100010";
        C <= "00010111";
        wait for clk_period;
        A <= "11010111";
        B <= "00011010";
        C <= "11000011";
        wait for clk_period;
        A <= "00011110";
        B <= "00000100";
        C <= "00011101";
        wait for clk_period;
        A <= "01001110";
        B <= "10110111";
        C <= "11010010";
        wait for clk_period;
        A <= "01010001";
        B <= "11111101";
        C <= "10000011";
        wait for clk_period;
        A <= "10010111";
        B <= "10111110";
        C <= "10111101";
        wait for clk_period;
        A <= "00111001";
        B <= "00111001";
        C <= "10011011";
        wait for clk_period;
        A <= "10001010";
        B <= "10111110";
        C <= "00010001";
        wait for clk_period;
        A <= "00000111";
        B <= "00111111";
        C <= "00110101";
        wait for clk_period;
        A <= "01110111";
        B <= "10001001";
        C <= "00111000";
        wait for clk_period;
        A <= "10111110";
        B <= "10100100";
        C <= "00110001";
        wait for clk_period;
        A <= "01101011";
        B <= "10101100";
        C <= "11101000";
        wait for clk_period;
        A <= "01110001";
        B <= "00001001";
        C <= "11000101";
        wait for clk_period;
        A <= "00011010";
        B <= "01010100";
        C <= "00110110";
        wait for clk_period;
        A <= "11100101";
        B <= "00010110";
        C <= "10101111";
        wait for clk_period;
        A <= "11011101";
        B <= "11000101";
        C <= "10111101";
        wait for clk_period;
        A <= "10111101";
        B <= "00001101";
        C <= "00101100";
        wait for clk_period;
        A <= "00101111";
        B <= "01000100";
        C <= "00100010";
        wait for clk_period;
        A <= "01110000";
        B <= "10100100";
        C <= "01100101";
        wait for clk_period;
        A <= "11100100";
        B <= "01111010";
        C <= "00010100";
        wait for clk_period;
        A <= "01100000";
        B <= "10111001";
        C <= "11111111";
        wait for clk_period;
        A <= "11110110";
        B <= "11011111";
        C <= "10110110";
        wait for clk_period;
        A <= "11101011";
        B <= "11100010";
        C <= "11111111";
        wait for clk_period;
        A <= "00000111";
        B <= "00000000";
        C <= "11011111";
        wait for clk_period;
        A <= "00010001";
        B <= "10011111";
        C <= "00010010";
        wait for clk_period;
        A <= "00111010";
        B <= "10010000";
        C <= "11100110";
        wait for clk_period;
        A <= "10101011";
        B <= "01010100";
        C <= "10000011";
        wait for clk_period;
        A <= "00110011";
        B <= "11101101";
        C <= "10101011";
        wait for clk_period;
        A <= "11000010";
        B <= "10010011";
        C <= "01111101";
        wait for clk_period;
        A <= "00001110";
        B <= "10110111";
        C <= "00010010";
        wait for clk_period;
        A <= "11000000";
        B <= "01001000";
        C <= "10100100";
        wait for clk_period;
        A <= "01011000";
        B <= "01101000";
        C <= "11100010";
        wait for clk_period;
        A <= "10100110";
        B <= "01010011";
        C <= "00011010";
        wait for clk_period;
        A <= "00010001";
        B <= "01110101";
        C <= "00010001";
        wait for clk_period;
        A <= "00100010";
        B <= "11001111";
        C <= "01010010";
        wait for clk_period;
        A <= "11011111";
        B <= "00111011";
        C <= "01111001";
        wait for clk_period;
        A <= "10010000";
        B <= "00111000";
        C <= "01011111";
        wait for clk_period;
        A <= "10111110";
        B <= "00001111";
        C <= "11011110";
        wait for clk_period;
        A <= "11101101";
        B <= "00010011";
        C <= "01100011";
        wait for clk_period;
        A <= "01101100";
        B <= "11110101";
        C <= "01010010";
        wait for clk_period;
        A <= "01110011";
        B <= "11101111";
        C <= "11000111";
        wait for clk_period;
        A <= "10100111";
        B <= "10001101";
        C <= "00110100";
        wait for clk_period;
        A <= "11011101";
        B <= "11001010";
        C <= "01011101";
        wait for clk_period;
        A <= "00011110";
        B <= "10011010";
        C <= "11101110";
        wait for clk_period;
        A <= "11110101";
        B <= "11100011";
        C <= "11100000";
        wait for clk_period;
        A <= "10001110";
        B <= "10110010";
        C <= "00011010";
        wait for clk_period;
        A <= "01110111";
        B <= "01011000";
        C <= "10110111";
        wait for clk_period;
        A <= "00011001";
        B <= "11011100";
        C <= "11010110";
        wait for clk_period;
        A <= "00111111";
        B <= "11101100";
        C <= "00000001";
        wait for clk_period;
        A <= "01101010";
        B <= "00010000";
        C <= "01100010";
        wait for clk_period;
        A <= "00100111";
        B <= "01001100";
        C <= "01111000";
        wait for clk_period;
        A <= "11100110";
        B <= "01001001";
        C <= "00000010";
        wait for clk_period;
        A <= "01000111";
        B <= "00010000";
        C <= "00111010";
        wait for clk_period;
        A <= "01000001";
        B <= "01001011";
        C <= "10101101";
        wait for clk_period;
        A <= "00010101";
        B <= "11011101";
        C <= "10001100";
        wait for clk_period;
        A <= "01101011";
        B <= "00010101";
        C <= "00001001";
        wait for clk_period;
        A <= "10110000";
        B <= "10101011";
        C <= "11000011";
        wait for clk_period;
        A <= "00110101";
        B <= "11000001";
        C <= "11110000";
        wait for clk_period;
        A <= "11011100";
        B <= "10111111";
        C <= "11011000";
        wait for clk_period;
        A <= "00010010";
        B <= "00001011";
        C <= "11000100";
        wait for clk_period;
        A <= "10110100";
        B <= "00001110";
        C <= "00000000";
        wait for clk_period;
        A <= "10011100";
        B <= "00110010";
        C <= "10010110";
        wait for clk_period;
        A <= "10011010";
        B <= "11010110";
        C <= "01110101";
        wait for clk_period;
        A <= "10001100";
        B <= "11010011";
        C <= "00000110";
        wait for clk_period;
        A <= "11010101";
        B <= "11100010";
        C <= "01000000";
        wait for clk_period;
        A <= "11011111";
        B <= "01011011";
        C <= "11110101";
        wait for clk_period;
        A <= "10111011";
        B <= "00011111";
        C <= "11101010";
        wait for clk_period;
        A <= "00100101";
        B <= "00001101";
        C <= "00001111";
        wait for clk_period;
        A <= "01010011";
        B <= "11111001";
        C <= "11110011";
        wait for clk_period;
        A <= "10001010";
        B <= "01000000";
        C <= "10010010";
        wait for clk_period;
        A <= "01100011";
        B <= "00101010";
        C <= "11100101";
        wait for clk_period;
        A <= "01100000";
        B <= "00111111";
        C <= "10110001";
        wait for clk_period;
        A <= "01110111";
        B <= "11011100";
        C <= "00110001";
        wait for clk_period;
        A <= "01011011";
        B <= "10101010";
        C <= "01011011";
        wait for clk_period;
        A <= "11101111";
        B <= "11010101";
        C <= "11010000";
        wait for clk_period;
        A <= "00011010";
        B <= "11011100";
        C <= "01111100";
        wait for clk_period;
        A <= "01101100";
        B <= "11101100";
        C <= "11111110";
        wait for clk_period;
        A <= "00000111";
        B <= "01100111";
        C <= "11110000";
        wait for clk_period;
        A <= "00100100";
        B <= "00011001";
        C <= "11101011";
        wait for clk_period;
        A <= "01011101";
        B <= "11101100";
        C <= "00100001";
        wait for clk_period;
        A <= "00101011";
        B <= "00011110";
        C <= "00011111";
        wait for clk_period;
        A <= "00110000";
        B <= "10100010";
        C <= "11010010";
        wait for clk_period;
        A <= "11100110";
        B <= "10101000";
        C <= "01101110";
        wait for clk_period;
        A <= "01111010";
        B <= "11101010";
        C <= "10101011";
        wait for clk_period;
        A <= "10100111";
        B <= "00010101";
        C <= "00101011";
        wait for clk_period;
        A <= "00110000";
        B <= "01100110";
        C <= "11111100";
        wait for clk_period;
        A <= "00100110";
        B <= "10111011";
        C <= "10100011";
        wait for clk_period;
        A <= "10000010";
        B <= "10100111";
        C <= "11110110";
        wait for clk_period;
        A <= "01011101";
        B <= "00101001";
        C <= "00010100";
        wait for clk_period;
        A <= "11100000";
        B <= "01110111";
        C <= "00000111";
        wait for clk_period;
        A <= "11010011";
        B <= "11100001";
        C <= "10111111";
        wait for clk_period;
        A <= "10111001";
        B <= "01011111";
        C <= "10100111";
        wait for clk_period;
        A <= "10001010";
        B <= "01000000";
        C <= "11101110";
        wait for clk_period;
        A <= "10101000";
        B <= "00010111";
        C <= "10110101";
        wait for clk_period;
        A <= "00011110";
        B <= "00101111";
        C <= "00011100";
        wait for clk_period;
        A <= "01011110";
        B <= "01010110";
        C <= "00001010";
        wait for clk_period;
        A <= "01011001";
        B <= "11111110";
        C <= "00001110";
        wait for clk_period;
        A <= "11110100";
        B <= "01010001";
        C <= "00001110";
        wait for clk_period;
        A <= "01111100";
        B <= "10011011";
        C <= "10101001";
        wait for clk_period;
        A <= "00011110";
        B <= "01001100";
        C <= "10111000";
        wait for clk_period;
        A <= "00110111";
        B <= "10100110";
        C <= "11100110";
        wait for clk_period;
        A <= "10011001";
        B <= "01011001";
        C <= "01101101";
        wait for clk_period;
        A <= "10100011";
        B <= "00111000";
        C <= "11101110";
        wait for clk_period;
        A <= "10101110";
        B <= "11011010";
        C <= "01111100";
        wait for clk_period;
        A <= "01011110";
        B <= "00000110";
        C <= "01111100";
        wait for clk_period;
        A <= "01010001";
        B <= "11011010";
        C <= "10110011";
        wait for clk_period;
        A <= "01001010";
        B <= "11110001";
        C <= "01100100";
        wait for clk_period;
        A <= "11100100";
        B <= "01010100";
        C <= "01100111";
        wait for clk_period;
        A <= "00111110";
        B <= "11010101";
        C <= "00111110";
        wait for clk_period;
        A <= "01101000";
        B <= "00101010";
        C <= "10010010";
        wait for clk_period;
        A <= "11101100";
        B <= "00110100";
        C <= "01101101";
        wait for clk_period;
        A <= "01001000";
        B <= "10101110";
        C <= "00010011";
        wait for clk_period;
        A <= "11011111";
        B <= "10111111";
        C <= "11110100";
        wait for clk_period;
        A <= "00111001";
        B <= "10000001";
        C <= "01101000";
        wait for clk_period;
        A <= "11010001";
        B <= "10110110";
        C <= "11111110";
        wait for clk_period;
        A <= "10110100";
        B <= "10111101";
        C <= "10111011";
        wait for clk_period;
        A <= "00101111";
        B <= "11000000";
        C <= "11110010";
        wait for clk_period;
        A <= "11010100";
        B <= "00001000";
        C <= "11010100";
        wait for clk_period;
        A <= "01011001";
        B <= "10111001";
        C <= "11101100";
        wait for clk_period;
        A <= "11010101";
        B <= "11100111";
        C <= "11101001";
        wait for clk_period;
        A <= "10010000";
        B <= "10111010";
        C <= "00100000";
        wait for clk_period;
        A <= "11101001";
        B <= "10110101";
        C <= "11111100";
        wait for clk_period;
        A <= "10101001";
        B <= "00111000";
        C <= "11100111";
        wait for clk_period;
        A <= "11100011";
        B <= "00001101";
        C <= "01100111";
        wait for clk_period;
        A <= "01011011";
        B <= "01111010";
        C <= "00110110";
        wait for clk_period;
        A <= "01111101";
        B <= "01010010";
        C <= "00001110";
        wait for clk_period;
        A <= "11110011";
        B <= "00001011";
        C <= "11110000";
        wait for clk_period;
        A <= "10110110";
        B <= "01110100";
        C <= "10000101";
        wait for clk_period;
        A <= "11110001";
        B <= "10101101";
        C <= "01110111";
        wait for clk_period;
        A <= "01000000";
        B <= "11100010";
        C <= "10010011";
        wait for clk_period;
        A <= "01000110";
        B <= "01001001";
        C <= "00110011";
        wait for clk_period;
        A <= "00100000";
        B <= "10001010";
        C <= "01101000";
        wait for clk_period;
        A <= "01110000";
        B <= "00101001";
        C <= "11111101";
        wait for clk_period;
        A <= "10011111";
        B <= "10011111";
        C <= "11110100";
        wait for clk_period;
        A <= "01000101";
        B <= "10001000";
        C <= "11111101";
        wait for clk_period;
        A <= "00100110";
        B <= "01000110";
        C <= "00100010";
        wait for clk_period;
        A <= "00010101";
        B <= "10000110";
        C <= "10111010";
        wait for clk_period;
        A <= "10110110";
        B <= "01111000";
        C <= "01000011";
        wait for clk_period;
        A <= "10001100";
        B <= "11111010";
        C <= "00101100";
        wait for clk_period;
        A <= "11001001";
        B <= "00000110";
        C <= "11011010";
        wait for clk_period;
        A <= "00101101";
        B <= "00000100";
        C <= "00010110";
        wait for clk_period;
        A <= "10110101";
        B <= "11011101";
        C <= "00010001";
        wait for clk_period;
        A <= "10101010";
        B <= "01001000";
        C <= "01100010";
        wait for clk_period;
        A <= "01100110";
        B <= "01100100";
        C <= "11101101";
        wait for clk_period;
        A <= "11000100";
        B <= "00110110";
        C <= "01100100";
        wait for clk_period;
        A <= "01101110";
        B <= "00111111";
        C <= "00000010";
        wait for clk_period;
        A <= "11000111";
        B <= "10001111";
        C <= "10011001";
        wait for clk_period;
        A <= "01011001";
        B <= "11101011";
        C <= "10000000";
        wait for clk_period;
        A <= "10100001";
        B <= "00100011";
        C <= "01011001";
        wait for clk_period;
        A <= "11110011";
        B <= "01010100";
        C <= "00001110";
        wait for clk_period;
        A <= "01111101";
        B <= "11000110";
        C <= "10110111";
        wait for clk_period;
        A <= "01110100";
        B <= "00111100";
        C <= "00110011";
        wait for clk_period;
        A <= "10011000";
        B <= "10001010";
        C <= "01011100";
        wait for clk_period;
        A <= "01001111";
        B <= "11011010";
        C <= "10001010";
        wait for clk_period;
        A <= "01011011";
        B <= "00101001";
        C <= "00011001";
        wait for clk_period;
        A <= "11111001";
        B <= "00111000";
        C <= "10101100";
        wait for clk_period;
        A <= "11101101";
        B <= "00010111";
        C <= "10110110";
        wait for clk_period;
        A <= "11000111";
        B <= "10100101";
        C <= "01100001";
        wait for clk_period;
        A <= "01011010";
        B <= "01011100";
        C <= "10011010";
        wait for clk_period;
        A <= "01100011";
        B <= "10010000";
        C <= "00001001";
        wait for clk_period;
        A <= "10111000";
        B <= "11011011";
        C <= "00110110";
        wait for clk_period;
        A <= "10110011";
        B <= "00111000";
        C <= "01000110";
        wait for clk_period;
        A <= "00010100";
        B <= "01001111";
        C <= "00001111";
        wait for clk_period;
        A <= "00000011";
        B <= "11010101";
        C <= "10010100";
        wait for clk_period;
        A <= "11100111";
        B <= "10101010";
        C <= "10111000";
        wait for clk_period;
        A <= "11101110";
        B <= "00000111";
        C <= "10011100";
        wait for clk_period;
        A <= "01100110";
        B <= "01011100";
        C <= "10001010";
        wait for clk_period;
        A <= "01001001";
        B <= "11101000";
        C <= "11010110";
        wait for clk_period;
        A <= "10010100";
        B <= "01100100";
        C <= "10111110";
        wait for clk_period;
        A <= "11111101";
        B <= "00100010";
        C <= "00001000";
        wait for clk_period;
        A <= "10101010";
        B <= "00111001";
        C <= "10010100";
        wait for clk_period;
        A <= "11110100";
        B <= "11110111";
        C <= "01001111";
        wait for clk_period;
        A <= "00110100";
        B <= "11011101";
        C <= "11010010";
        wait for clk_period;
        A <= "11110001";
        B <= "10001001";
        C <= "01010000";
        wait for clk_period;
        A <= "11101010";
        B <= "00000000";
        C <= "10111100";
        wait for clk_period;
        A <= "10011100";
        B <= "01100101";
        C <= "10100011";
        wait for clk_period;
        A <= "00000100";
        B <= "11111001";
        C <= "11110001";
        wait for clk_period;
        A <= "01111111";
        B <= "10011101";
        C <= "00011111";
        wait for clk_period;
        A <= "11011101";
        B <= "01110111";
        C <= "10010001";
        wait for clk_period;
        A <= "01111011";
        B <= "10011100";
        C <= "00100011";
        wait for clk_period;
        A <= "01000111";
        B <= "01111111";
        C <= "10001010";
        wait for clk_period;
        A <= "00001101";
        B <= "10101000";
        C <= "00110011";
        wait for clk_period;
        A <= "01100100";
        B <= "10100100";
        C <= "01011001";
        wait for clk_period;
        A <= "10101100";
        B <= "11011100";
        C <= "00011011";
        wait for clk_period;
        A <= "10110111";
        B <= "00011000";
        C <= "01100011";
        wait for clk_period;
        A <= "10000100";
        B <= "10011011";
        C <= "00000100";
        wait for clk_period;
        A <= "10111101";
        B <= "11110011";
        C <= "10000111";
        wait for clk_period;
        A <= "11101000";
        B <= "00000100";
        C <= "11110001";
        wait for clk_period;
        A <= "00001001";
        B <= "11111011";
        C <= "01001101";
        wait for clk_period;
        A <= "11110000";
        B <= "00011100";
        C <= "10111101";
        wait for clk_period;
        A <= "01001010";
        B <= "01010110";
        C <= "10011011";
        wait for clk_period;
        A <= "01101011";
        B <= "01011100";
        C <= "01001001";
        wait for clk_period;
        A <= "00110111";
        B <= "01011110";
        C <= "00110001";
        wait for clk_period;
        A <= "10100101";
        B <= "01001010";
        C <= "11111110";
        wait for clk_period;
        A <= "10100101";
        B <= "10101010";
        C <= "00001010";
        wait for clk_period;
        A <= "01010111";
        B <= "01110111";
        C <= "00111110";
        wait for clk_period;
        A <= "01110001";
        B <= "11000101";
        C <= "10011001";
        wait for clk_period;
        A <= "01010010";
        B <= "00101111";
        C <= "01111011";
        wait for clk_period;
        A <= "01001000";
        B <= "10001010";
        C <= "00000100";
        wait for clk_period;
        A <= "00110111";
        B <= "01001111";
        C <= "10010001";
        wait for clk_period;
        A <= "10001001";
        B <= "11001000";
        C <= "10100010";
        wait for clk_period;
        A <= "10101000";
        B <= "01010001";
        C <= "11111011";
        wait for clk_period;
        A <= "01010010";
        B <= "10101000";
        C <= "10011001";
        wait for clk_period;
        A <= "00000010";
        B <= "01000111";
        C <= "10101001";
        wait for clk_period;
        A <= "01101101";
        B <= "01100100";
        C <= "00100101";
        wait for clk_period;
        A <= "11000010";
        B <= "11110110";
        C <= "10000110";
        wait for clk_period;
        A <= "10011100";
        B <= "10111111";
        C <= "11001001";
        wait for clk_period;
        A <= "00110001";
        B <= "10000110";
        C <= "01011111";
        wait for clk_period;
        A <= "11110001";
        B <= "11101111";
        C <= "01010011";
        wait for clk_period;
        A <= "11010001";
        B <= "11001100";
        C <= "00110101";
        wait for clk_period;
        A <= "01101001";
        B <= "01011010";
        C <= "00110110";
        wait for clk_period;
        A <= "10000001";
        B <= "01010000";
        C <= "01101000";
        wait for clk_period;
        A <= "01000011";
        B <= "10000111";
        C <= "00110110";
        wait for clk_period;
        A <= "11100001";
        B <= "11010111";
        C <= "11011001";
        wait for clk_period;
        A <= "10111100";
        B <= "11010000";
        C <= "10100100";
        wait for clk_period;
        A <= "11011010";
        B <= "00001100";
        C <= "00011010";
        wait for clk_period;
        A <= "10101100";
        B <= "00110001";
        C <= "00010110";
        wait for clk_period;
        A <= "10100011";
        B <= "00101000";
        C <= "11110110";
        wait for clk_period;
        A <= "00010011";
        B <= "10100111";
        C <= "10011001";
        wait for clk_period;
        A <= "11001011";
        B <= "10010100";
        C <= "10101110";
        wait for clk_period;
        A <= "01001100";
        B <= "00111111";
        C <= "11111100";
        wait for clk_period;
        A <= "11101011";
        B <= "11001111";
        C <= "11010011";
        wait for clk_period;
        A <= "10100110";
        B <= "01100001";
        C <= "10110101";
        wait for clk_period;
        A <= "10011001";
        B <= "11100110";
        C <= "11101001";
        wait for clk_period;
        A <= "01110011";
        B <= "10010110";
        C <= "10001000";
        wait for clk_period;
        A <= "10100010";
        B <= "00000000";
        C <= "00110001";
        wait for clk_period;
        A <= "11100010";
        B <= "00101111";
        C <= "01110001";
        wait for clk_period;
        A <= "11011100";
        B <= "10011100";
        C <= "10110001";
        wait for clk_period;
        A <= "00001110";
        B <= "11100100";
        C <= "10101001";
        wait for clk_period;
        A <= "10001000";
        B <= "10001111";
        C <= "00110001";
        wait for clk_period;
        A <= "00100101";
        B <= "11011110";
        C <= "11000101";
        wait for clk_period;
        A <= "01101101";
        B <= "11001100";
        C <= "10100110";
        wait for clk_period;
        A <= "11001111";
        B <= "11001100";
        C <= "01010000";
        wait for clk_period;
        A <= "11001000";
        B <= "01011111";
        C <= "11101011";
        wait for clk_period;
        A <= "10111000";
        B <= "01111000";
        C <= "10111111";
        wait for clk_period;
        A <= "00000111";
        B <= "10110010";
        C <= "00111101";
        wait for clk_period;
        A <= "01110100";
        B <= "01001011";
        C <= "10100100";
        wait for clk_period;
        A <= "00001011";
        B <= "01001001";
        C <= "10010001";
        wait for clk_period;
        A <= "11010100";
        B <= "11000110";
        C <= "11010000";
        wait for clk_period;
        A <= "10110111";
        B <= "11100111";
        C <= "00010110";
        wait for clk_period;
        A <= "00110011";
        B <= "10111000";
        C <= "10101001";
        wait for clk_period;
        A <= "10001011";
        B <= "00001101";
        C <= "10110111";
        wait for clk_period;
        A <= "10011100";
        B <= "01101001";
        C <= "10011000";
        wait for clk_period;
        A <= "01010000";
        B <= "10101011";
        C <= "00111011";
        wait for clk_period;
        A <= "01001010";
        B <= "11100101";
        C <= "00011000";
        wait for clk_period;
        A <= "10011100";
        B <= "00100000";
        C <= "10010101";
        wait for clk_period;
        A <= "10011011";
        B <= "01010000";
        C <= "00001000";
        wait for clk_period;
        A <= "00110000";
        B <= "01000110";
        C <= "10010100";
        wait for clk_period;
        A <= "10100110";
        B <= "00101001";
        C <= "10010101";
        wait for clk_period;
        A <= "10010001";
        B <= "00000111";
        C <= "01001101";
        wait for clk_period;
        A <= "01011101";
        B <= "10111101";
        C <= "01010010";
        wait for clk_period;
        A <= "11010111";
        B <= "00000100";
        C <= "11101101";
        wait for clk_period;
        A <= "11010011";
        B <= "11101110";
        C <= "10001001";
        wait for clk_period;
        A <= "10001000";
        B <= "11000100";
        C <= "11010101";
        wait for clk_period;
        A <= "01001000";
        B <= "11111110";
        C <= "01111011";
        wait for clk_period;
        A <= "11010011";
        B <= "01111011";
        C <= "10001001";
        wait for clk_period;
        A <= "11000000";
        B <= "01101011";
        C <= "10101011";
        wait for clk_period;
        A <= "00100011";
        B <= "01100100";
        C <= "00000000";
        wait for clk_period;
        A <= "10011100";
        B <= "01011010";
        C <= "11000011";
        wait for clk_period;
        A <= "10111000";
        B <= "10011100";
        C <= "01101011";
        wait for clk_period;
        A <= "01011110";
        B <= "00010101";
        C <= "11010010";
        wait for clk_period;
        A <= "11100001";
        B <= "11110011";
        C <= "10101111";
        wait for clk_period;
        A <= "11100110";
        B <= "00110010";
        C <= "11011001";
        wait for clk_period;
        A <= "01011011";
        B <= "01000000";
        C <= "10000101";
        wait for clk_period;
        A <= "10000100";
        B <= "00010110";
        C <= "00010001";
        wait for clk_period;
        A <= "10000010";
        B <= "00100011";
        C <= "11000110";
        wait for clk_period;
        A <= "01001010";
        B <= "11101011";
        C <= "00100100";
        wait for clk_period;
        A <= "01100000";
        B <= "01010010";
        C <= "10100110";
        wait for clk_period;
        A <= "01011000";
        B <= "00110101";
        C <= "00100110";
        wait for clk_period;
        A <= "00000110";
        B <= "10110110";
        C <= "10110111";
        wait for clk_period;
        A <= "00111101";
        B <= "10100011";
        C <= "11110111";
        wait for clk_period;
        A <= "00111110";
        B <= "11101101";
        C <= "01101101";
        wait for clk_period;
        A <= "10110011";
        B <= "00111110";
        C <= "00111100";
        wait for clk_period;
        A <= "01000111";
        B <= "11100011";
        C <= "00010111";
        wait for clk_period;
        A <= "10000010";
        B <= "10010110";
        C <= "00010000";
        wait for clk_period;
        A <= "10010110";
        B <= "01111011";
        C <= "10011110";
        wait for clk_period;
        A <= "10101001";
        B <= "11010011";
        C <= "11011011";
        wait for clk_period;
        A <= "00001000";
        B <= "00100010";
        C <= "10111100";
        wait for clk_period;
        A <= "01110010";
        B <= "10011111";
        C <= "01101000";
        wait for clk_period;
        A <= "11000110";
        B <= "10010010";
        C <= "01101011";
        wait for clk_period;
        A <= "10010100";
        B <= "01111100";
        C <= "10010001";
        wait for clk_period;
        A <= "01110100";
        B <= "01101111";
        C <= "11110000";
        wait for clk_period;
        A <= "11111011";
        B <= "01011010";
        C <= "10110011";
        wait for clk_period;
        A <= "00100101";
        B <= "11001010";
        C <= "01101111";
        wait for clk_period;
        A <= "11101101";
        B <= "10000011";
        C <= "10101001";
        wait for clk_period;
        A <= "10100001";
        B <= "10011000";
        C <= "01001001";
        wait for clk_period;
        A <= "10110010";
        B <= "01011011";
        C <= "11110010";
        wait for clk_period;
        A <= "00101100";
        B <= "01010010";
        C <= "10011010";
        wait for clk_period;
        A <= "01101001";
        B <= "01001000";
        C <= "10110010";
        wait for clk_period;
        A <= "00010011";
        B <= "00011100";
        C <= "11011000";
        wait for clk_period;
        A <= "11100101";
        B <= "01110110";
        C <= "00101001";
        wait for clk_period;
        A <= "10001001";
        B <= "10101100";
        C <= "01110101";
        wait for clk_period;
        A <= "00011100";
        B <= "11000001";
        C <= "01011011";
        wait for clk_period;
        A <= "10011101";
        B <= "11111100";
        C <= "01010111";
        wait for clk_period;
        A <= "11101010";
        B <= "00110001";
        C <= "00110111";
        wait for clk_period;
        A <= "00001000";
        B <= "11111110";
        C <= "11010100";
        wait for clk_period;
        A <= "01110011";
        B <= "01010011";
        C <= "00011011";
        wait for clk_period;
        A <= "11001000";
        B <= "00110110";
        C <= "00000001";
        wait for clk_period;
        A <= "00001011";
        B <= "01000101";
        C <= "11001100";
        wait for clk_period;
        A <= "00011111";
        B <= "10001101";
        C <= "11011100";
        wait for clk_period;
        A <= "00000000";
        B <= "00010110";
        C <= "00111101";
        wait for clk_period;
        A <= "00100010";
        B <= "00000011";
        C <= "01111110";
        wait for clk_period;
        A <= "00110100";
        B <= "01011100";
        C <= "10001111";
        wait for clk_period;
        A <= "01100011";
        B <= "01110010";
        C <= "01110101";
        wait for clk_period;
        A <= "01000010";
        B <= "10101101";
        C <= "01001010";
        wait for clk_period;
        A <= "01111110";
        B <= "11101110";
        C <= "01000100";
        wait for clk_period;
        A <= "11000110";
        B <= "01111011";
        C <= "11001001";
        wait for clk_period;
        A <= "00100100";
        B <= "10010000";
        C <= "11100111";
        wait for clk_period;
        A <= "11001000";
        B <= "11001101";
        C <= "11111011";
        wait for clk_period;
        A <= "00110001";
        B <= "00111001";
        C <= "01011110";
        wait for clk_period;
        A <= "11000111";
        B <= "00111001";
        C <= "00100010";
        wait for clk_period;
        A <= "11100010";
        B <= "11001001";
        C <= "11011001";
        wait for clk_period;
        A <= "01111011";
        B <= "01101110";
        C <= "01110010";
        wait for clk_period;
        A <= "10011100";
        B <= "01011111";
        C <= "11001010";
        wait for clk_period;
        A <= "01110110";
        B <= "00100100";
        C <= "00001111";
        wait for clk_period;
        A <= "10110000";
        B <= "10110010";
        C <= "00100111";
        wait for clk_period;
        A <= "11000110";
        B <= "00000111";
        C <= "10111100";
        wait for clk_period;
        A <= "10101111";
        B <= "10110001";
        C <= "11001011";
        wait for clk_period;
        A <= "11101110";
        B <= "11110000";
        C <= "11000001";
        wait for clk_period;
        A <= "01000110";
        B <= "01010011";
        C <= "00001111";
        wait for clk_period;
        A <= "10100000";
        B <= "11000110";
        C <= "01010100";
        wait for clk_period;
        A <= "10110001";
        B <= "00000000";
        C <= "10000100";
        wait for clk_period;
        A <= "10001001";
        B <= "11001000";
        C <= "01110010";
        wait for clk_period;
        A <= "01000111";
        B <= "10011000";
        C <= "00100001";
        wait for clk_period;
        A <= "10100000";
        B <= "01101101";
        C <= "11011011";
        wait for clk_period;
        A <= "00111000";
        B <= "10111101";
        C <= "11111111";
        wait for clk_period;
        A <= "00101010";
        B <= "10100011";
        C <= "11100010";
        wait for clk_period;
        A <= "01110011";
        B <= "01001101";
        C <= "10101000";
        wait for clk_period;
        A <= "01110001";
        B <= "11011110";
        C <= "10111110";
        wait for clk_period;
        A <= "00011011";
        B <= "00011100";
        C <= "00110010";
        wait for clk_period;
        A <= "01101000";
        B <= "01100000";
        C <= "10100011";
        wait for clk_period;
        A <= "10101100";
        B <= "01000000";
        C <= "10010101";
        wait for clk_period;
        A <= "01010100";
        B <= "10100000";
        C <= "10011010";
        wait for clk_period;
        A <= "10010101";
        B <= "01110001";
        C <= "11000110";
        wait for clk_period;
        A <= "00100101";
        B <= "00001010";
        C <= "10100001";
        wait for clk_period;
        A <= "11011010";
        B <= "00010011";
        C <= "01110101";
        wait for clk_period;
        A <= "00100000";
        B <= "11011011";
        C <= "11100100";
        wait for clk_period;
        A <= "11110111";
        B <= "10110100";
        C <= "10111001";
        wait for clk_period;
        A <= "10000111";
        B <= "00001111";
        C <= "10110100";
        wait for clk_period;
        A <= "00100110";
        B <= "01111100";
        C <= "01010011";
        wait for clk_period;
        A <= "10010011";
        B <= "11001100";
        C <= "01010100";
        wait for clk_period;
        A <= "11010001";
        B <= "01101000";
        C <= "00100010";
        wait for clk_period;
        A <= "11110100";
        B <= "01000101";
        C <= "10000010";
        wait for clk_period;
        A <= "10000110";
        B <= "10011110";
        C <= "11111011";
        wait for clk_period;
        A <= "00100100";
        B <= "11000010";
        C <= "01011101";
        wait for clk_period;
        A <= "10101100";
        B <= "11100110";
        C <= "01010011";
        wait for clk_period;
        A <= "10111111";
        B <= "01110001";
        C <= "10100110";
        wait for clk_period;
        A <= "01000111";
        B <= "11110001";
        C <= "10001100";
        wait for clk_period;
        A <= "10101010";
        B <= "11111100";
        C <= "01100111";
        wait for clk_period;
        A <= "10101001";
        B <= "00001100";
        C <= "10011100";
        wait for clk_period;
        A <= "01010110";
        B <= "00011001";
        C <= "00000000";
        wait for clk_period;
        A <= "11000010";
        B <= "01111011";
        C <= "01010011";
        wait for clk_period;
        A <= "00110110";
        B <= "11000011";
        C <= "10011010";
        wait for clk_period;
        A <= "00111011";
        B <= "01001101";
        C <= "00101110";
        wait for clk_period;
        A <= "01000110";
        B <= "01001111";
        C <= "10000110";
        wait for clk_period;
        A <= "10010000";
        B <= "01000100";
        C <= "11000101";
        wait for clk_period;
        A <= "11101111";
        B <= "00011011";
        C <= "10010110";
        wait for clk_period;
        A <= "01010101";
        B <= "01010110";
        C <= "00001101";
        wait for clk_period;
        A <= "01011010";
        B <= "00101001";
        C <= "00011001";
        wait for clk_period;
        A <= "00110000";
        B <= "10000001";
        C <= "11110000";
        wait for clk_period;
        A <= "00011010";
        B <= "00111101";
        C <= "01100000";
        wait for clk_period;
        A <= "01101111";
        B <= "10000100";
        C <= "11000101";
        wait for clk_period;
        A <= "10000010";
        B <= "01101101";
        C <= "00000001";
        wait for clk_period;
        A <= "10110111";
        B <= "10111011";
        C <= "00001101";
        wait for clk_period;
        A <= "10101100";
        B <= "00011010";
        C <= "11010010";
        wait for clk_period;
        A <= "01010001";
        B <= "00111001";
        C <= "11000011";
        wait for clk_period;
        A <= "01001011";
        B <= "11101011";
        C <= "00011000";
        wait for clk_period;
        A <= "11001100";
        B <= "11010000";
        C <= "01100110";
        wait for clk_period;
        A <= "11110110";
        B <= "01010101";
        C <= "00000000";
        wait for clk_period;
        A <= "01010100";
        B <= "01111110";
        C <= "10001010";
        wait for clk_period;
        A <= "01011001";
        B <= "10100000";
        C <= "11110011";
        wait for clk_period;
        A <= "10000101";
        B <= "00010010";
        C <= "00011010";
        wait for clk_period;
        A <= "01011011";
        B <= "00111100";
        C <= "10110011";
        wait for clk_period;
        A <= "00100110";
        B <= "10111101";
        C <= "10111010";
        wait for clk_period;
        A <= "01000011";
        B <= "00100011";
        C <= "00110100";
        wait for clk_period;
        A <= "10111101";
        B <= "11000011";
        C <= "11000000";
        wait for clk_period;
        A <= "01000000";
        B <= "11011011";
        C <= "11111101";
        wait for clk_period;
        A <= "01111100";
        B <= "10111110";
        C <= "00011001";
        wait for clk_period;
        A <= "01011111";
        B <= "01101111";
        C <= "10110101";
        wait for clk_period;
        A <= "10101000";
        B <= "01100011";
        C <= "00001011";
        wait for clk_period;
        A <= "11101001";
        B <= "11001000";
        C <= "01001101";
        wait for clk_period;
        A <= "10010000";
        B <= "10110111";
        C <= "10001101";
        wait for clk_period;
        A <= "00101011";
        B <= "11111100";
        C <= "01100010";
        wait for clk_period;
        A <= "10111101";
        B <= "11101101";
        C <= "10111111";
        wait for clk_period;
        A <= "11011001";
        B <= "00000110";
        C <= "10101011";
        wait for clk_period;
        A <= "00101110";
        B <= "01010000";
        C <= "10010010";
        wait for clk_period;
        A <= "01100101";
        B <= "00110100";
        C <= "11110110";
        wait for clk_period;
        A <= "00111111";
        B <= "01110000";
        C <= "11000011";
        wait for clk_period;
        A <= "10111010";
        B <= "10101101";
        C <= "00110000";
        wait for clk_period;
        A <= "00010101";
        B <= "11101110";
        C <= "10010001";
        wait for clk_period;
        A <= "01100011";
        B <= "11100010";
        C <= "01101110";
        wait for clk_period;
        A <= "11100101";
        B <= "11010011";
        C <= "10011010";
        wait for clk_period;
        A <= "00000110";
        B <= "01011001";
        C <= "10000101";
        wait for clk_period;
        A <= "11010001";
        B <= "00000110";
        C <= "01001100";
        wait for clk_period;
        A <= "10011110";
        B <= "10011101";
        C <= "00001111";
        wait for clk_period;
        A <= "01011111";
        B <= "11011001";
        C <= "01100011";
        wait for clk_period;
        A <= "00101111";
        B <= "10101010";
        C <= "00001110";
        wait for clk_period;
        A <= "11000010";
        B <= "00000111";
        C <= "01110001";
        wait for clk_period;
        A <= "00111011";
        B <= "10001010";
        C <= "00000100";
        wait for clk_period;
        A <= "01001000";
        B <= "10001110";
        C <= "10010001";
        wait for clk_period;
        A <= "00101111";
        B <= "11000100";
        C <= "10011111";
        wait for clk_period;
        A <= "10100101";
        B <= "10000110";
        C <= "00000100";
        wait for clk_period;
        A <= "01001110";
        B <= "10111101";
        C <= "01011010";
        wait for clk_period;
        A <= "11000100";
        B <= "11011111";
        C <= "10001111";
        wait for clk_period;
        A <= "11100111";
        B <= "11101100";
        C <= "11001000";
        wait for clk_period;
        A <= "11011001";
        B <= "00001110";
        C <= "11101100";
        wait for clk_period;
        A <= "01101110";
        B <= "10100111";
        C <= "10011011";
        wait for clk_period;
        A <= "00100010";
        B <= "11001101";
        C <= "00100110";
        wait for clk_period;
        A <= "10010111";
        B <= "10101110";
        C <= "11111110";
        wait for clk_period;
        A <= "10110110";
        B <= "10111101";
        C <= "00111101";
        wait for clk_period;
        A <= "10011110";
        B <= "11111001";
        C <= "00000001";
        wait for clk_period;
        A <= "01011100";
        B <= "00101100";
        C <= "01100010";
        wait for clk_period;
        A <= "00111101";
        B <= "01001000";
        C <= "10100100";
        wait for clk_period;
        A <= "01011010";
        B <= "10001110";
        C <= "10010110";
        wait for clk_period;
        A <= "11101111";
        B <= "11111101";
        C <= "00101011";
        wait for clk_period;
        A <= "11111010";
        B <= "01100010";
        C <= "10001010";
        wait for clk_period;
        A <= "00101100";
        B <= "01111100";
        C <= "10011011";
        wait for clk_period;
        A <= "00110110";
        B <= "00110000";
        C <= "00100101";
        wait for clk_period;
        A <= "11001010";
        B <= "01110111";
        C <= "10011011";
        wait for clk_period;
        A <= "10010110";
        B <= "11010001";
        C <= "11101100";
        wait for clk_period;
        A <= "11101000";
        B <= "11101110";
        C <= "00100110";
        wait for clk_period;
        A <= "00101001";
        B <= "00100101";
        C <= "10100011";
        wait for clk_period;
        A <= "11011111";
        B <= "00010110";
        C <= "01000000";
        wait for clk_period;
        A <= "01001110";
        B <= "00001011";
        C <= "01111010";
        wait for clk_period;
        A <= "11110010";
        B <= "10011101";
        C <= "01001100";
        wait for clk_period;
        A <= "01110000";
        B <= "01001110";
        C <= "11011101";
        wait for clk_period;
        A <= "10011111";
        B <= "01011000";
        C <= "11110001";
        wait for clk_period;
        A <= "00101000";
        B <= "10010011";
        C <= "10010100";
        wait for clk_period;
        A <= "10101001";
        B <= "10110110";
        C <= "11111000";
        wait for clk_period;
        A <= "10111111";
        B <= "11100011";
        C <= "10010011";
        wait for clk_period;
        A <= "01001011";
        B <= "11100000";
        C <= "01000010";
        wait for clk_period;
        A <= "10111000";
        B <= "11110100";
        C <= "10100100";
        wait for clk_period;
        A <= "01101010";
        B <= "00001010";
        C <= "10110000";
        wait for clk_period;
        A <= "10011100";
        B <= "11000000";
        C <= "00011101";
        wait for clk_period;
        A <= "01101010";
        B <= "10001110";
        C <= "00100101";
        wait for clk_period;
        A <= "01001001";
        B <= "11011011";
        C <= "01001001";
        wait for clk_period;
        A <= "01001001";
        B <= "11111011";
        C <= "11000010";
        wait for clk_period;
        A <= "10101000";
        B <= "11110000";
        C <= "00101100";
        wait for clk_period;
        A <= "10010110";
        B <= "01001001";
        C <= "10100100";
        wait for clk_period;
        A <= "10000100";
        B <= "00001010";
        C <= "10110110";
        wait for clk_period;
        A <= "01000001";
        B <= "10011001";
        C <= "01101010";
        wait for clk_period;
        A <= "10001100";
        B <= "00001110";
        C <= "10000110";
        wait for clk_period;
        A <= "10110011";
        B <= "10001100";
        C <= "10101010";
        wait for clk_period;
        A <= "01111110";
        B <= "01110101";
        C <= "10101011";
        wait for clk_period;
        A <= "00010111";
        B <= "11100000";
        C <= "10110000";
        wait for clk_period;
        A <= "11000101";
        B <= "10001001";
        C <= "10100100";
        wait for clk_period;
        A <= "01001110";
        B <= "11011100";
        C <= "00110001";
        wait for clk_period;
        A <= "10110101";
        B <= "01101111";
        C <= "10110101";
        wait for clk_period;
        A <= "10110000";
        B <= "11110101";
        C <= "11010101";
        wait for clk_period;
        A <= "00110000";
        B <= "00110100";
        C <= "11101110";
        wait for clk_period;
        A <= "00000110";
        B <= "01100110";
        C <= "10011011";
        wait for clk_period;
        A <= "01111100";
        B <= "00111000";
        C <= "10110101";
        wait for clk_period;
        A <= "01011001";
        B <= "11110110";
        C <= "01000101";
        wait for clk_period;
        A <= "11100001";
        B <= "11010000";
        C <= "10101001";
        wait for clk_period;
        A <= "01010010";
        B <= "10001001";
        C <= "00010000";
        wait for clk_period;
        A <= "00101011";
        B <= "00001000";
        C <= "01101101";
        wait for clk_period;
        A <= "00111110";
        B <= "01111001";
        C <= "11001111";
        wait for clk_period;
        A <= "00010010";
        B <= "00111001";
        C <= "10000010";
        wait for clk_period;
        A <= "11100001";
        B <= "10111000";
        C <= "11011001";
        wait for clk_period;
        A <= "11000010";
        B <= "00010011";
        C <= "01000100";
        wait for clk_period;
        A <= "00011001";
        B <= "11100111";
        C <= "11000001";
        wait for clk_period;
        A <= "10000110";
        B <= "01101101";
        C <= "11011010";
        wait for clk_period;
        A <= "11101001";
        B <= "00110011";
        C <= "01011010";
        wait for clk_period;
        A <= "11011101";
        B <= "00010111";
        C <= "11001001";
        wait for clk_period;
        A <= "11110001";
        B <= "00011001";
        C <= "10001110";
        wait for clk_period;
        A <= "11000010";
        B <= "11010101";
        C <= "10001101";
        wait for clk_period;
        A <= "10100001";
        B <= "10001010";
        C <= "01001100";
        wait for clk_period;
        A <= "11100110";
        B <= "11100101";
        C <= "10101100";
        wait for clk_period;
        A <= "11111010";
        B <= "01010100";
        C <= "01110000";
        wait for clk_period;
        A <= "10110110";
        B <= "01000000";
        C <= "01010000";
        wait for clk_period;
        A <= "11000010";
        B <= "11000010";
        C <= "00111011";
        wait for clk_period;
        A <= "10000000";
        B <= "01001100";
        C <= "00011000";
        wait for clk_period;
        A <= "11000011";
        B <= "01010110";
        C <= "11100010";
        wait for clk_period;
        A <= "11000011";
        B <= "11101110";
        C <= "00101111";
        wait for clk_period;
        A <= "11100111";
        B <= "11000000";
        C <= "00010111";
        wait for clk_period;
        A <= "01101111";
        B <= "00100001";
        C <= "10110011";
        wait for clk_period;
        A <= "01101001";
        B <= "01011001";
        C <= "00111000";
        wait for clk_period;
        A <= "11001111";
        B <= "00011010";
        C <= "01000010";
        wait for clk_period;
        A <= "00111100";
        B <= "10000111";
        C <= "01100011";
        wait for clk_period;
        A <= "01111001";
        B <= "01101111";
        C <= "00011001";
        wait for clk_period;
        A <= "10011111";
        B <= "10010111";
        C <= "11100111";
        wait for clk_period;
        A <= "00100110";
        B <= "01010111";
        C <= "00011101";
        wait for clk_period;
        A <= "11110101";
        B <= "00100001";
        C <= "11001001";
        wait for clk_period;
        A <= "01101011";
        B <= "01001000";
        C <= "10101100";
        wait for clk_period;
        A <= "11011001";
        B <= "00000001";
        C <= "10101010";
        wait for clk_period;
        A <= "11110001";
        B <= "11010011";
        C <= "01110010";
        wait for clk_period;
        A <= "01110101";
        B <= "01100000";
        C <= "00101000";
        wait for clk_period;
        A <= "10101101";
        B <= "00111001";
        C <= "10001100";
        wait for clk_period;
        A <= "01111000";
        B <= "11001101";
        C <= "01111110";
        wait for clk_period;
        A <= "01111110";
        B <= "11101001";
        C <= "10111011";
        wait for clk_period;
        A <= "00101100";
        B <= "00010110";
        C <= "00011010";
        wait for clk_period;
        A <= "10011111";
        B <= "01011000";
        C <= "10111100";
        wait for clk_period;
        A <= "00110000";
        B <= "01111000";
        C <= "00001100";
        wait for clk_period;
        A <= "01010101";
        B <= "10101011";
        C <= "10000001";
        wait for clk_period;
        A <= "11110110";
        B <= "10111101";
        C <= "11011001";
        wait for clk_period;
        A <= "01110101";
        B <= "10110000";
        C <= "10110110";
        wait for clk_period;
        A <= "00111110";
        B <= "11011111";
        C <= "00110101";
        wait for clk_period;
        A <= "10110110";
        B <= "00010101";
        C <= "01110111";
        wait for clk_period;
        A <= "10001000";
        B <= "01110000";
        C <= "00110111";
        wait for clk_period;
        A <= "11000100";
        B <= "01000110";
        C <= "10011000";
        wait for clk_period;
        A <= "11110111";
        B <= "10010001";
        C <= "00100000";
        wait for clk_period;
        A <= "10111000";
        B <= "10011100";
        C <= "00101000";
        wait for clk_period;
        A <= "00111111";
        B <= "11101110";
        C <= "01000101";
        wait for clk_period;
        A <= "11110000";
        B <= "00101010";
        C <= "01101101";
        wait for clk_period;
        A <= "10011001";
        B <= "10001100";
        C <= "00001110";
        wait for clk_period;
        A <= "10111111";
        B <= "10011011";
        C <= "00110110";
        wait for clk_period;
        A <= "01001110";
        B <= "10000000";
        C <= "00100101";
        wait for clk_period;
        A <= "11100001";
        B <= "00110011";
        C <= "10111101";
        wait for clk_period;
        A <= "01100110";
        B <= "01010011";
        C <= "11010100";
        wait for clk_period;
        A <= "10000100";
        B <= "11111101";
        C <= "11110011";
        wait for clk_period;
        A <= "01001010";
        B <= "00010101";
        C <= "01101101";
        wait for clk_period;
        A <= "01101010";
        B <= "01001001";
        C <= "01010100";
        wait for clk_period;
        A <= "11000110";
        B <= "10000111";
        C <= "00001100";
        wait for clk_period;
        A <= "01101100";
        B <= "10001100";
        C <= "01101100";
        wait for clk_period;
        A <= "01010010";
        B <= "11110011";
        C <= "11001010";
        wait for clk_period;
        A <= "01011100";
        B <= "00110011";
        C <= "11100000";
        wait for clk_period;
        A <= "11111101";
        B <= "00100000";
        C <= "01011110";
        wait for clk_period;
        A <= "01001010";
        B <= "01110000";
        C <= "01110001";
        wait for clk_period;
        A <= "00110010";
        B <= "10100000";
        C <= "11001101";
        wait for clk_period;
        A <= "10001111";
        B <= "10101110";
        C <= "01010010";
        wait for clk_period;
        A <= "00101000";
        B <= "11011111";
        C <= "10011011";
        wait for clk_period;
        A <= "11100001";
        B <= "11110001";
        C <= "11011100";
        wait for clk_period;
        A <= "11100110";
        B <= "11100101";
        C <= "10111001";
        wait for clk_period;
        A <= "11000101";
        B <= "11110010";
        C <= "00110000";
        wait for clk_period;
        A <= "11011000";
        B <= "11011000";
        C <= "00010101";
        wait for clk_period;
        A <= "00101101";
        B <= "11110000";
        C <= "00110100";
        wait for clk_period;
        A <= "00111011";
        B <= "01101111";
        C <= "01000010";
        wait for clk_period;
        A <= "11111000";
        B <= "11011111";
        C <= "00100000";
        wait for clk_period;
        A <= "00010011";
        B <= "00111100";
        C <= "10010001";
        wait for clk_period;
        A <= "10110100";
        B <= "00010001";
        C <= "01010001";
        wait for clk_period;
        A <= "01110010";
        B <= "10010101";
        C <= "00101001";
        wait for clk_period;
        A <= "11001101";
        B <= "11001100";
        C <= "01111001";
        wait for clk_period;
        A <= "11010000";
        B <= "00111101";
        C <= "10010110";
        wait for clk_period;
        A <= "00111001";
        B <= "01101111";
        C <= "10100011";
        wait for clk_period;
        A <= "00000011";
        B <= "11100101";
        C <= "11010101";
        wait for clk_period;
        A <= "00111110";
        B <= "11111100";
        C <= "10101101";
        wait for clk_period;
        A <= "00111111";
        B <= "11010100";
        C <= "00100010";
        wait for clk_period;
        A <= "01101001";
        B <= "01000100";
        C <= "11101000";
        wait for clk_period;
        A <= "11111010";
        B <= "10110010";
        C <= "00010110";
        wait for clk_period;
        A <= "11011100";
        B <= "01011011";
        C <= "10000000";
        wait for clk_period;
        A <= "10011001";
        B <= "11110000";
        C <= "01111011";
        wait for clk_period;
        A <= "10001110";
        B <= "01111000";
        C <= "00000010";
        wait for clk_period;
        A <= "00010011";
        B <= "00001100";
        C <= "10110011";
        wait for clk_period;
        A <= "00100111";
        B <= "11110111";
        C <= "00111111";
        wait for clk_period;
        A <= "01101100";
        B <= "11000111";
        C <= "10010011";
        wait for clk_period;
        A <= "10111101";
        B <= "11100001";
        C <= "11011111";
        wait for clk_period;
        A <= "00000010";
        B <= "01010010";
        C <= "11111111";
        wait for clk_period;
        A <= "01010101";
        B <= "01111101";
        C <= "10010110";
        wait for clk_period;
        A <= "01001101";
        B <= "00000110";
        C <= "10101010";
        wait for clk_period;
        A <= "00000101";
        B <= "01101110";
        C <= "00101111";
        wait for clk_period;
        A <= "01000101";
        B <= "01001101";
        C <= "01011000";
        wait for clk_period;
        A <= "01001011";
        B <= "01000000";
        C <= "00110101";
        wait for clk_period;
        A <= "11100100";
        B <= "01110101";
        C <= "00111011";
        wait for clk_period;
        A <= "00010101";
        B <= "10111111";
        C <= "00111001";
        wait for clk_period;
        A <= "10011011";
        B <= "10100111";
        C <= "01001101";
        wait for clk_period;
        A <= "00001010";
        B <= "10101010";
        C <= "11001010";
        wait for clk_period;
        A <= "01000000";
        B <= "11011110";
        C <= "10011110";
        wait for clk_period;
        A <= "10001000";
        B <= "00111111";
        C <= "11001110";
        wait for clk_period;
        A <= "11010110";
        B <= "11001101";
        C <= "10111010";
        wait for clk_period;
        A <= "00001110";
        B <= "00101101";
        C <= "01110101";
        wait for clk_period;
        A <= "10101010";
        B <= "01000001";
        C <= "01010010";
        wait for clk_period;
        A <= "10110110";
        B <= "11001101";
        C <= "01101110";
        wait for clk_period;
        A <= "01010101";
        B <= "00000000";
        C <= "00010010";
        wait for clk_period;
        A <= "01110011";
        B <= "11011110";
        C <= "01010100";
        wait for clk_period;
        A <= "01011101";
        B <= "10111110";
        C <= "00011100";
        wait for clk_period;
        A <= "10000001";
        B <= "00100101";
        C <= "11001001";
        wait for clk_period;
        A <= "01110000";
        B <= "01001110";
        C <= "11101010";
        wait for clk_period;
        A <= "00010101";
        B <= "01011001";
        C <= "10001110";
        wait for clk_period;
        A <= "00100110";
        B <= "00110100";
        C <= "00010111";
        wait for clk_period;
        A <= "00110010";
        B <= "01111100";
        C <= "11101000";
        wait for clk_period;
        A <= "01111110";
        B <= "00000101";
        C <= "11001001";
        wait for clk_period;
        A <= "11001010";
        B <= "10110001";
        C <= "10001010";
        wait for clk_period;
        A <= "10011001";
        B <= "00100100";
        C <= "10111010";
        wait for clk_period;
        A <= "00101100";
        B <= "00101100";
        C <= "11000101";
        wait for clk_period;
        A <= "10010001";
        B <= "10010111";
        C <= "10010111";
        wait for clk_period;
        A <= "11101100";
        B <= "10010101";
        C <= "11000101";
        wait for clk_period;
        A <= "01111000";
        B <= "10101011";
        C <= "11100000";
        wait for clk_period;
        A <= "00101010";
        B <= "11000011";
        C <= "11011100";
        wait for clk_period;
        A <= "00001010";
        B <= "11100010";
        C <= "00001111";
        wait for clk_period;
        A <= "01000000";
        B <= "10100011";
        C <= "10110110";
        wait for clk_period;
        A <= "01111110";
        B <= "10000110";
        C <= "10100000";
        wait for clk_period;
        A <= "10010111";
        B <= "11011000";
        C <= "00010111";
        wait for clk_period;
        A <= "10010011";
        B <= "01100101";
        C <= "10111000";
        wait for clk_period;
        A <= "00110101";
        B <= "10100100";
        C <= "11011010";
        wait for clk_period;
        A <= "01010011";
        B <= "10001011";
        C <= "01010101";
        wait for clk_period;
        A <= "11110101";
        B <= "01101110";
        C <= "01111001";
        wait for clk_period;
        A <= "11100110";
        B <= "01110101";
        C <= "00000011";
        wait for clk_period;
        A <= "01111101";
        B <= "10001000";
        C <= "10010101";
        wait for clk_period;
        A <= "00010011";
        B <= "11100000";
        C <= "01011110";
        wait for clk_period;
        A <= "00110010";
        B <= "00110100";
        C <= "00110110";
        wait for clk_period;
        A <= "01110110";
        B <= "01111111";
        C <= "10101111";
        wait for clk_period;
        A <= "00100111";
        B <= "10111101";
        C <= "01011000";
        wait for clk_period;
        A <= "11001001";
        B <= "10011110";
        C <= "00000110";
        wait for clk_period;
        A <= "11010110";
        B <= "10001010";
        C <= "00101110";
        wait for clk_period;
        A <= "11110011";
        B <= "10001110";
        C <= "11100010";
        wait for clk_period;
        A <= "10110011";
        B <= "01001100";
        C <= "10011110";
        wait for clk_period;
        A <= "01010111";
        B <= "00010001";
        C <= "01010111";
        wait for clk_period;
        A <= "11100011";
        B <= "10011000";
        C <= "01100101";
        wait for clk_period;
        A <= "10000100";
        B <= "00111000";
        C <= "00001011";
        wait for clk_period;
        A <= "01111111";
        B <= "00101010";
        C <= "10010000";
        wait for clk_period;
        A <= "00010110";
        B <= "11000100";
        C <= "01100010";
        wait for clk_period;
        A <= "11111010";
        B <= "11100100";
        C <= "11011110";
        wait for clk_period;
        A <= "11111101";
        B <= "01101110";
        C <= "10010000";
        wait for clk_period;
        A <= "11100110";
        B <= "10001011";
        C <= "10100111";
        wait for clk_period;
        A <= "11100011";
        B <= "11011110";
        C <= "01001001";
        wait for clk_period;
        A <= "01001101";
        B <= "11011000";
        C <= "00010000";
        wait for clk_period;
        A <= "10101111";
        B <= "11110001";
        C <= "00000001";
        wait for clk_period;
        A <= "01011100";
        B <= "11101101";
        C <= "11110001";
        wait for clk_period;
        A <= "00111011";
        B <= "11000000";
        C <= "01101011";
        wait for clk_period;
        A <= "11101101";
        B <= "00000110";
        C <= "01001010";
        wait for clk_period;
        A <= "01011111";
        B <= "00101011";
        C <= "01001100";
        wait for clk_period;
        A <= "01110001";
        B <= "01011101";
        C <= "11110111";
        wait for clk_period;
        A <= "00111000";
        B <= "11010010";
        C <= "00010001";
        wait for clk_period;
        A <= "10010110";
        B <= "00010110";
        C <= "00101111";
        wait for clk_period;
        A <= "11110011";
        B <= "10101101";
        C <= "00010000";
        wait for clk_period;
        A <= "10100011";
        B <= "10101111";
        C <= "10100110";
        wait for clk_period;
        A <= "11001000";
        B <= "00010110";
        C <= "00101110";
        wait for clk_period;
        A <= "11110010";
        B <= "10101111";
        C <= "01111010";
        wait for clk_period;
        A <= "10110100";
        B <= "10010111";
        C <= "11011100";
        wait for clk_period;
        A <= "00011001";
        B <= "11000000";
        C <= "11110000";
        wait for clk_period;
        A <= "10110111";
        B <= "01100101";
        C <= "00011111";
        wait for clk_period;
        A <= "10001000";
        B <= "01001000";
        C <= "01001001";
        wait for clk_period;
        A <= "00001001";
        B <= "10110011";
        C <= "00010111";
        wait for clk_period;
        A <= "11101011";
        B <= "01100000";
        C <= "01111001";
        wait for clk_period;
        A <= "11110111";
        B <= "01011111";
        C <= "00110000";
        wait for clk_period;
        A <= "00100101";
        B <= "10000010";
        C <= "11111001";
        wait for clk_period;
        A <= "10001100";
        B <= "00011110";
        C <= "00010101";
        wait for clk_period;
        A <= "00100011";
        B <= "01100111";
        C <= "01010000";
        wait for clk_period;
        A <= "11111000";
        B <= "10001101";
        C <= "01011010";
        wait for clk_period;
        A <= "11001000";
        B <= "11010001";
        C <= "10000010";
        wait for clk_period;
        A <= "00110110";
        B <= "01001011";
        C <= "10001101";
        wait for clk_period;
        A <= "00100001";
        B <= "11010011";
        C <= "00100100";
        wait for clk_period;
        A <= "11111000";
        B <= "11011000";
        C <= "10101000";
        wait for clk_period;
        A <= "10000000";
        B <= "01100101";
        C <= "01111000";
        wait for clk_period;
        A <= "10000010";
        B <= "10101100";
        C <= "10000001";
        wait for clk_period;
        A <= "00001010";
        B <= "00100011";
        C <= "11010111";
        wait for clk_period;
        A <= "00001011";
        B <= "11110010";
        C <= "00010110";
        wait for clk_period;
        A <= "11101011";
        B <= "10011001";
        C <= "10101110";
        wait for clk_period;
        A <= "01011101";
        B <= "00010000";
        C <= "00001101";
        wait for clk_period;
        A <= "01010010";
        B <= "01110011";
        C <= "01011111";
        wait for clk_period;
        A <= "00111111";
        B <= "11101000";
        C <= "01000100";
        wait for clk_period;
        A <= "11100100";
        B <= "11110111";
        C <= "01010000";
        wait for clk_period;
        A <= "10010001";
        B <= "01000110";
        C <= "01100100";
        wait for clk_period;
        A <= "00110111";
        B <= "01010000";
        C <= "11100100";
        wait for clk_period;
        A <= "10111111";
        B <= "10000111";
        C <= "10101111";
        wait for clk_period;
        A <= "00100110";
        B <= "11011101";
        C <= "11010001";
        wait for clk_period;
        A <= "00011000";
        B <= "01000111";
        C <= "11010000";
        wait for clk_period;
        A <= "11011100";
        B <= "01010110";
        C <= "00111111";
        wait for clk_period;
        A <= "11111100";
        B <= "01100011";
        C <= "00010011";
        wait for clk_period;
        A <= "01001101";
        B <= "11111011";
        C <= "10101100";
        wait for clk_period;
        A <= "00010110";
        B <= "11010100";
        C <= "10001010";
        wait for clk_period;
        A <= "11001010";
        B <= "00101100";
        C <= "01010000";
        wait for clk_period;
        A <= "00001011";
        B <= "10001101";
        C <= "11011011";
        wait for clk_period;
        A <= "01111000";
        B <= "10010001";
        C <= "10100110";
        wait for clk_period;
        A <= "00000111";
        B <= "01100101";
        C <= "01101101";
        wait for clk_period;
        A <= "10011011";
        B <= "10011010";
        C <= "10010100";
        wait for clk_period;
        A <= "01000101";
        B <= "11100100";
        C <= "11100000";
        wait for clk_period;
        A <= "10011011";
        B <= "11101110";
        C <= "10100000";
        wait for clk_period;
        A <= "11011111";
        B <= "11101101";
        C <= "10111010";
        wait for clk_period;
        A <= "10000000";
        B <= "11110011";
        C <= "00100010";
        wait for clk_period;
        A <= "01010001";
        B <= "11101110";
        C <= "00101010";
        wait for clk_period;
        A <= "00111111";
        B <= "10101001";
        C <= "10000100";
        wait for clk_period;
        A <= "11110101";
        B <= "11110000";
        C <= "01000101";
        wait for clk_period;
        A <= "11111011";
        B <= "10101110";
        C <= "00100011";
        wait for clk_period;
        A <= "10000111";
        B <= "10101010";
        C <= "00001110";
        wait for clk_period;
        A <= "11111111";
        B <= "11110011";
        C <= "11110000";
        wait for clk_period;
        A <= "00011111";
        B <= "10000111";
        C <= "10100011";
        wait for clk_period;
        A <= "01100001";
        B <= "11110000";
        C <= "10001011";
        wait for clk_period;
        A <= "01010000";
        B <= "01101011";
        C <= "10001011";
        wait for clk_period;
        A <= "11111001";
        B <= "10100010";
        C <= "11100011";
        wait for clk_period;
        A <= "01001010";
        B <= "10011011";
        C <= "10101111";
        wait for clk_period;
        A <= "10001001";
        B <= "01111101";
        C <= "01000100";
        wait for clk_period;
        A <= "01011010";
        B <= "10010111";
        C <= "01101110";
        wait for clk_period;
        A <= "11011111";
        B <= "11001011";
        C <= "00100110";
        wait for clk_period;
        A <= "01000101";
        B <= "01000001";
        C <= "10000100";
        wait for clk_period;
        A <= "10001111";
        B <= "00100010";
        C <= "01111100";
        wait for clk_period;
        A <= "11110110";
        B <= "01100011";
        C <= "00000100";
        wait for clk_period;
        A <= "11010011";
        B <= "10010001";
        C <= "01100111";
        wait for clk_period;
        A <= "01011010";
        B <= "11011010";
        C <= "10101111";
        wait for clk_period;
        A <= "00110001";
        B <= "01011111";
        C <= "10011011";
        wait for clk_period;
        A <= "00110110";
        B <= "11100001";
        C <= "01110000";
        wait for clk_period;
        A <= "11001100";
        B <= "01011111";
        C <= "10101101";
        wait for clk_period;
        A <= "11010000";
        B <= "01111110";
        C <= "00111010";
        wait for clk_period;
        A <= "10100100";
        B <= "11010011";
        C <= "11110111";
        wait for clk_period;
        A <= "01011001";
        B <= "00101001";
        C <= "11100110";
        wait for clk_period;
        A <= "00101110";
        B <= "11001101";
        C <= "11110001";
        wait for clk_period;
        A <= "11000011";
        B <= "11101100";
        C <= "00001110";
        wait for clk_period;
        A <= "10010000";
        B <= "00101100";
        C <= "00111111";
        wait for clk_period;
        A <= "10101010";
        B <= "00110010";
        C <= "01101100";
        wait for clk_period;
        A <= "10101110";
        B <= "00100001";
        C <= "00101111";
        wait for clk_period;
        A <= "11010011";
        B <= "11101000";
        C <= "01011101";
        wait for clk_period;
        A <= "11010101";
        B <= "10010010";
        C <= "01011001";
        wait for clk_period;
        A <= "10001111";
        B <= "11010100";
        C <= "01000010";
        wait for clk_period;
        A <= "00110100";
        B <= "00110100";
        C <= "00001001";
        wait for clk_period;
        A <= "10000111";
        B <= "00100100";
        C <= "00001011";
        wait for clk_period;
        A <= "11001111";
        B <= "11011101";
        C <= "10111111";
        wait for clk_period;
        A <= "10111110";
        B <= "10101111";
        C <= "01001001";
        wait for clk_period;
        A <= "00110001";
        B <= "10000110";
        C <= "10101100";
        wait for clk_period;
        A <= "01100110";
        B <= "01000110";
        C <= "01001001";
        wait for clk_period;
        A <= "10001101";
        B <= "00000010";
        C <= "10001010";
        wait for clk_period;
        A <= "00011000";
        B <= "10000100";
        C <= "10011000";
        wait for clk_period;
        A <= "10110100";
        B <= "10010011";
        C <= "01100111";
        wait for clk_period;
        A <= "10000000";
        B <= "11111100";
        C <= "10011011";
        wait for clk_period;
        A <= "00011110";
        B <= "00000001";
        C <= "11100101";
        wait for clk_period;
        A <= "00011111";
        B <= "10011101";
        C <= "11011101";
        wait for clk_period;
        A <= "11110011";
        B <= "01110111";
        C <= "10101100";
        wait for clk_period;
        A <= "10100111";
        B <= "00100001";
        C <= "11110011";
        wait for clk_period;
        A <= "01111010";
        B <= "01110001";
        C <= "01100001";
        wait for clk_period;
        A <= "00011111";
        B <= "00101000";
        C <= "01100001";
        wait for clk_period;
        A <= "11110010";
        B <= "01111110";
        C <= "11100110";
        wait for clk_period;
        A <= "01001010";
        B <= "10010110";
        C <= "00001111";
        wait for clk_period;
        A <= "11001110";
        B <= "11000110";
        C <= "11101011";
        wait for clk_period;
        A <= "11111011";
        B <= "00100101";
        C <= "11100001";
        wait for clk_period;
        A <= "00011010";
        B <= "01101100";
        C <= "10101000";
        wait for clk_period;
        A <= "11001000";
        B <= "01101100";
        C <= "01110001";
        wait for clk_period;
        A <= "11100011";
        B <= "10010000";
        C <= "10101010";
        wait for clk_period;
        A <= "00100011";
        B <= "10101101";
        C <= "10010101";
        wait for clk_period;
        A <= "10100111";
        B <= "00011111";
        C <= "10000111";
        wait for clk_period;
        A <= "00001100";
        B <= "11001100";
        C <= "01011101";
        wait for clk_period;
        A <= "10101001";
        B <= "01110011";
        C <= "00011110";
        wait for clk_period;
        A <= "01110000";
        B <= "00010111";
        C <= "11100100";
        wait for clk_period;
        A <= "00111001";
        B <= "10010001";
        C <= "10101101";
        wait for clk_period;
        A <= "11100111";
        B <= "11111011";
        C <= "11111000";
        wait for clk_period;
        A <= "10000000";
        B <= "11111111";
        C <= "11001011";
        wait for clk_period;
        A <= "11001100";
        B <= "01101000";
        C <= "00001011";
        wait for clk_period;
        A <= "11101110";
        B <= "00101110";
        C <= "11110110";
        wait for clk_period;
        A <= "01110111";
        B <= "01110111";
        C <= "10010100";
        wait for clk_period;
        A <= "10110001";
        B <= "00011101";
        C <= "11111111";
        wait for clk_period;
        A <= "01001011";
        B <= "01010101";
        C <= "01101011";
        wait for clk_period;
        A <= "01110101";
        B <= "11110011";
        C <= "11010010";
        wait for clk_period;
        A <= "01000100";
        B <= "01000000";
        C <= "11010110";
        wait for clk_period;
        A <= "00110111";
        B <= "00100010";
        C <= "10011000";
        wait for clk_period;
        A <= "00010101";
        B <= "10000001";
        C <= "11111001";
        wait for clk_period;
        A <= "11011101";
        B <= "01010010";
        C <= "10111011";
        wait for clk_period;
        A <= "01110110";
        B <= "11101111";
        C <= "00011011";
        wait for clk_period;
        A <= "11000010";
        B <= "11111001";
        C <= "11101010";
        wait for clk_period;
        A <= "11001000";
        B <= "11110101";
        C <= "00100001";
        wait for clk_period;
        A <= "01010001";
        B <= "00111100";
        C <= "00010000";
        wait for clk_period;
        A <= "11111111";
        B <= "11101111";
        C <= "00110001";
        wait for clk_period;
        A <= "11101011";
        B <= "11100111";
        C <= "01010010";
        wait for clk_period;
        A <= "11011011";
        B <= "11001000";
        C <= "10000111";
        wait for clk_period;
        A <= "11100111";
        B <= "01000010";
        C <= "00001001";
        wait for clk_period;
        A <= "00101011";
        B <= "11100001";
        C <= "10110011";
        wait for clk_period;
        A <= "11111100";
        B <= "10001101";
        C <= "01000011";
        wait for clk_period;
        A <= "00101100";
        B <= "00010011";
        C <= "10100010";
        wait for clk_period;
        A <= "11000001";
        B <= "11000111";
        C <= "01101111";
        wait for clk_period;
        A <= "00111010";
        B <= "10110001";
        C <= "01011111";
        wait for clk_period;
        A <= "00000110";
        B <= "11010010";
        C <= "10011100";
        wait for clk_period;
        A <= "11001010";
        B <= "10011101";
        C <= "01110101";
        wait for clk_period;
        A <= "11100001";
        B <= "01100100";
        C <= "01101110";
        wait for clk_period;
        A <= "01001101";
        B <= "01000000";
        C <= "00010011";
        wait for clk_period;
        A <= "10100110";
        B <= "01110000";
        C <= "10110101";
        wait for clk_period;
        A <= "11000011";
        B <= "01111010";
        C <= "11010010";
        wait for clk_period;
        A <= "11010101";
        B <= "00011111";
        C <= "01011011";
        wait for clk_period;
        A <= "00100100";
        B <= "01011010";
        C <= "01011110";
        wait for clk_period;
        A <= "00001110";
        B <= "11001110";
        C <= "00110110";
        wait for clk_period;
        A <= "10001111";
        B <= "11011110";
        C <= "11101000";
        wait for clk_period;
        A <= "01100100";
        B <= "11010000";
        C <= "10110100";
        wait for clk_period;
        A <= "01011011";
        B <= "11001100";
        C <= "11011111";
        wait for clk_period;
        A <= "10010111";
        B <= "00110000";
        C <= "00110101";
        wait for clk_period;
        A <= "01101110";
        B <= "01110001";
        C <= "01111010";
        wait for clk_period;
        A <= "00001011";
        B <= "00101001";
        C <= "00101100";
        wait for clk_period;
        A <= "00011101";
        B <= "11111000";
        C <= "00110101";
        wait for clk_period;
        A <= "01100101";
        B <= "11001100";
        C <= "11110111";
        wait for clk_period;
        A <= "00100000";
        B <= "00100001";
        C <= "00110000";
        wait for clk_period;
        A <= "10101110";
        B <= "01010111";
        C <= "00110010";
        wait for clk_period;
        A <= "01101111";
        B <= "10110000";
        C <= "10110000";
        wait for clk_period;
        A <= "11001000";
        B <= "01000101";
        C <= "11110101";
        wait for clk_period;
        A <= "01010010";
        B <= "00100001";
        C <= "11000111";
        wait for clk_period;
        A <= "10100101";
        B <= "00110000";
        C <= "11010001";
        wait for clk_period;
        A <= "01111100";
        B <= "11110001";
        C <= "11101001";
        wait for clk_period;
        A <= "01111100";
        B <= "10110011";
        C <= "01011111";
        wait for clk_period;
        A <= "11000101";
        B <= "11010100";
        C <= "10100100";
        wait for clk_period;
        A <= "11101011";
        B <= "11010110";
        C <= "00010011";
        wait for clk_period;
        A <= "11011001";
        B <= "11011011";
        C <= "01011111";
        wait for clk_period;
        A <= "01111001";
        B <= "01000111";
        C <= "00010110";
        wait for clk_period;
        A <= "11001100";
        B <= "00111111";
        C <= "11101010";
        wait for clk_period;
        A <= "11010111";
        B <= "11111101";
        C <= "01011100";
        wait for clk_period;
        A <= "11001101";
        B <= "00000011";
        C <= "01000101";
        wait for clk_period;
        A <= "00001001";
        B <= "11000110";
        C <= "10110011";
        wait for clk_period;
        A <= "11101000";
        B <= "11000000";
        C <= "10011111";
        wait for clk_period;
        A <= "00111101";
        B <= "01010110";
        C <= "10011111";
        wait for clk_period;
        A <= "11111101";
        B <= "00010010";
        C <= "10111110";
        wait for clk_period;
        A <= "10111001";
        B <= "01100111";
        C <= "11000011";
        wait for clk_period;
        A <= "01100111";
        B <= "00110111";
        C <= "10001101";
        wait for clk_period;
        A <= "01000101";
        B <= "01111011";
        C <= "10010111";
        wait for clk_period;
        A <= "00100100";
        B <= "11001111";
        C <= "01011011";
        wait for clk_period;
        A <= "10111001";
        B <= "10111001";
        C <= "01000110";
        wait for clk_period;
        A <= "11011111";
        B <= "11011001";
        C <= "00101000";
        wait for clk_period;
        A <= "11000110";
        B <= "01000011";
        C <= "10011001";
        wait for clk_period;
        A <= "11010001";
        B <= "10000011";
        C <= "01101111";
        wait for clk_period;
        A <= "11100000";
        B <= "01100000";
        C <= "00010001";
        wait for clk_period;
        A <= "01000011";
        B <= "00100110";
        C <= "11001011";
        wait for clk_period;
        A <= "01010001";
        B <= "00011000";
        C <= "01001100";
        wait for clk_period;
        A <= "01000010";
        B <= "00010101";
        C <= "00101011";
        wait for clk_period;
        A <= "11110000";
        B <= "01000101";
        C <= "01101111";
        wait for clk_period;
        A <= "11100010";
        B <= "01111011";
        C <= "01000111";
        wait for clk_period;
        A <= "10000000";
        B <= "11010010";
        C <= "00100010";
        wait for clk_period;
        A <= "11100110";
        B <= "11101110";
        C <= "10001110";
        wait for clk_period;
        A <= "01011110";
        B <= "10111110";
        C <= "10111111";
        wait for clk_period;
        A <= "00100000";
        B <= "01101111";
        C <= "00010010";
        wait for clk_period;
        A <= "00100101";
        B <= "00010101";
        C <= "10100010";
        wait for clk_period;
        A <= "11100000";
        B <= "00011110";
        C <= "10101000";
        wait for clk_period;
        A <= "10100111";
        B <= "01100010";
        C <= "00111101";
        wait for clk_period;
        A <= "00101001";
        B <= "11001001";
        C <= "10110100";
        wait for clk_period;
        A <= "00001000";
        B <= "00101101";
        C <= "01011010";
        wait for clk_period;
        A <= "00101101";
        B <= "11010111";
        C <= "11011101";
        wait for clk_period;
        A <= "00101110";
        B <= "11010101";
        C <= "01010001";
        wait for clk_period;
        A <= "11111101";
        B <= "11100011";
        C <= "10110010";
        wait for clk_period;
        A <= "10010000";
        B <= "01010000";
        C <= "10001100";
        wait for clk_period;
        A <= "11011001";
        B <= "01110110";
        C <= "10011111";
        wait for clk_period;
        A <= "11000001";
        B <= "01011110";
        C <= "00101110";
        wait for clk_period;
        A <= "11000110";
        B <= "11011001";
        C <= "01000011";
        wait for clk_period;
        A <= "11000011";
        B <= "00001000";
        C <= "11101110";
        wait for clk_period;
        A <= "11001100";
        B <= "11100101";
        C <= "10101001";
        wait for clk_period;
        A <= "11101010";
        B <= "01011001";
        C <= "10001110";
        wait for clk_period;
        A <= "01100110";
        B <= "10101101";
        C <= "01000111";
        wait for clk_period;
        A <= "10111100";
        B <= "00000101";
        C <= "10000110";
        wait for clk_period;
        A <= "01010000";
        B <= "00110000";
        C <= "10110011";
        wait for clk_period;
        A <= "00110110";
        B <= "00000100";
        C <= "01100001";
        wait for clk_period;
        A <= "10101110";
        B <= "11010000";
        C <= "00010100";
        wait for clk_period;
        A <= "11011001";
        B <= "11011100";
        C <= "10010011";
        wait for clk_period;
        A <= "11111011";
        B <= "00011111";
        C <= "11110110";
        wait for clk_period;
        A <= "11000101";
        B <= "01001101";
        C <= "10001111";
        wait for clk_period;
        A <= "00001000";
        B <= "01101100";
        C <= "01111001";
        wait for clk_period;
        A <= "11110111";
        B <= "00010000";
        C <= "01000000";
        wait for clk_period;
        A <= "00001111";
        B <= "11011111";
        C <= "00100101";
        wait for clk_period;
        A <= "01101010";
        B <= "00111001";
        C <= "11111010";
        wait for clk_period;
        A <= "10011010";
        B <= "11100110";
        C <= "10001111";
        wait for clk_period;
        A <= "10101101";
        B <= "00111000";
        C <= "11011100";
        wait for clk_period;
        A <= "10010101";
        B <= "00010111";
        C <= "01000111";
        wait for clk_period;
        A <= "00011101";
        B <= "11111011";
        C <= "00001000";
        wait for clk_period;
        A <= "00001100";
        B <= "10100111";
        C <= "11000100";
        wait for clk_period;
        A <= "10101100";
        B <= "00000011";
        C <= "00010101";
        wait for clk_period;
        A <= "11001000";
        B <= "01011100";
        C <= "11011110";
        wait for clk_period;
        A <= "10011000";
        B <= "01111100";
        C <= "00101100";
        wait for clk_period;
        A <= "10000101";
        B <= "10011000";
        C <= "11001001";
        wait for clk_period;
        A <= "11010110";
        B <= "10101100";
        C <= "11010110";
        wait for clk_period;
        A <= "11111010";
        B <= "11100101";
        C <= "00111010";
        wait for clk_period;
        A <= "10110100";
        B <= "10101111";
        C <= "11010010";
        wait for clk_period;
        A <= "01111110";
        B <= "01110010";
        C <= "10011101";
        wait for clk_period;
        A <= "11001000";
        B <= "01111011";
        C <= "10111000";
        wait for clk_period;
        A <= "10011101";
        B <= "01011011";
        C <= "11111100";
        wait for clk_period;
        A <= "11010001";
        B <= "10100011";
        C <= "01101001";
        wait for clk_period;
        A <= "10111000";
        B <= "10001110";
        C <= "10110100";
        wait for clk_period;
        A <= "01111110";
        B <= "11111111";
        C <= "00001111";
        wait for clk_period;
        A <= "00111101";
        B <= "10001101";
        C <= "01001111";
        wait for clk_period;
        A <= "01100000";
        B <= "10100010";
        C <= "11010111";
        wait for clk_period;
        A <= "01000111";
        B <= "00110001";
        C <= "01101111";
        wait for clk_period;
        A <= "01110110";
        B <= "01101010";
        C <= "00101100";
        wait for clk_period;
        A <= "01001011";
        B <= "10011100";
        C <= "01010111";
        wait for clk_period;
        A <= "00001011";
        B <= "00101111";
        C <= "01111100";
        wait for clk_period;
        A <= "00001101";
        B <= "10010001";
        C <= "10110010";
        wait for clk_period;
        A <= "01101011";
        B <= "11011110";
        C <= "00001110";
        wait for clk_period;
        A <= "10110000";
        B <= "11001001";
        C <= "11010010";
        wait for clk_period;
        A <= "10101101";
        B <= "00100001";
        C <= "10111011";
        wait for clk_period;
        A <= "01111100";
        B <= "01111110";
        C <= "10100100";
        wait for clk_period;
        A <= "11100000";
        B <= "00100001";
        C <= "01110001";
        wait for clk_period;
        A <= "10010110";
        B <= "01001000";
        C <= "11100010";
        wait for clk_period;
        A <= "00100100";
        B <= "01010110";
        C <= "00111000";
        wait for clk_period;
        A <= "11000101";
        B <= "00010001";
        C <= "10010001";
        wait for clk_period;
        A <= "11000100";
        B <= "10001100";
        C <= "10110111";
        wait for clk_period;
        A <= "10100101";
        B <= "10000101";
        C <= "11010101";
        wait for clk_period;
        A <= "10100101";
        B <= "11110000";
        C <= "11011000";
        wait for clk_period;
        A <= "01100000";
        B <= "11101000";
        C <= "11101100";
        wait for clk_period;
        A <= "11100001";
        B <= "10110100";
        C <= "01100010";
        wait for clk_period;
        A <= "11000000";
        B <= "01000011";
        C <= "01001110";
        wait for clk_period;
        A <= "00001110";
        B <= "01111101";
        C <= "10100100";
        wait for clk_period;
        A <= "00100010";
        B <= "10101011";
        C <= "01100101";
        wait for clk_period;
        A <= "10100001";
        B <= "01010111";
        C <= "10000100";
        wait for clk_period;
        A <= "01111101";
        B <= "11100100";
        C <= "10110101";
        wait for clk_period;
        A <= "00001101";
        B <= "10110101";
        C <= "01001011";
        wait for clk_period;
        A <= "11011111";
        B <= "00001001";
        C <= "10011100";
        wait for clk_period;
        A <= "01011001";
        B <= "01100001";
        C <= "00010000";
        wait for clk_period;
        A <= "11111010";
        B <= "00110011";
        C <= "00000100";
        wait for clk_period;
        A <= "10111100";
        B <= "00000100";
        C <= "11000101";
        wait for clk_period;
        A <= "11101001";
        B <= "00011111";
        C <= "00000000";
        wait for clk_period;
        A <= "01010010";
        B <= "10011001";
        C <= "11101011";
        wait for clk_period;
        A <= "10010100";
        B <= "00101011";
        C <= "11000111";
        wait for clk_period;
        A <= "00001101";
        B <= "10001101";
        C <= "00110101";
        wait for clk_period;
        A <= "01111000";
        B <= "00011000";
        C <= "00010001";
        wait for clk_period;
        A <= "01111101";
        B <= "01100000";
        C <= "00101010";
        wait for clk_period;
        A <= "00011000";
        B <= "01101101";
        C <= "11111110";
        wait for clk_period;
        A <= "10110110";
        B <= "10110000";
        C <= "00001001";
        wait for clk_period;
        A <= "00011100";
        B <= "00011001";
        C <= "10100101";
        wait for clk_period;
        A <= "00100000";
        B <= "10011110";
        C <= "11101010";
        wait for clk_period;
        A <= "10000010";
        B <= "01101001";
        C <= "11000011";
        wait for clk_period;
        A <= "11000011";
        B <= "01011000";
        C <= "10001001";
        wait for clk_period;
        A <= "10011011";
        B <= "01000010";
        C <= "11000001";
        wait for clk_period;
        A <= "01100101";
        B <= "10000000";
        C <= "11010110";
        wait for clk_period;
        A <= "00001101";
        B <= "00111010";
        C <= "00100011";
        wait for clk_period;
        A <= "01110001";
        B <= "10011100";
        C <= "01011011";
        wait for clk_period;
        A <= "01110000";
        B <= "00000110";
        C <= "00001110";
        wait for clk_period;
        A <= "10100100";
        B <= "00101010";
        C <= "11001101";
        wait for clk_period;
        A <= "10000011";
        B <= "00000000";
        C <= "01011000";
        wait for clk_period;
        A <= "11111011";
        B <= "10100010";
        C <= "00001001";
        wait for clk_period;
        A <= "11010100";
        B <= "10001000";
        C <= "10001000";
        wait for clk_period;
        A <= "10001100";
        B <= "01100011";
        C <= "11100011";
        wait for clk_period;
        A <= "00111001";
        B <= "11101011";
        C <= "00110111";
        wait for clk_period;
        A <= "11001110";
        B <= "11111011";
        C <= "10100100";
        wait for clk_period;
        A <= "11111111";
        B <= "01110000";
        C <= "00011110";
        wait for clk_period;
        A <= "01100110";
        B <= "00101011";
        C <= "11100010";
        wait for clk_period;
        A <= "10111110";
        B <= "00110101";
        C <= "00110011";
        wait for clk_period;
        A <= "11101011";
        B <= "00101010";
        C <= "00111001";
        wait for clk_period;
        A <= "11101110";
        B <= "11010001";
        C <= "00001001";
        wait for clk_period;
        A <= "00010011";
        B <= "11111100";
        C <= "01110001";
        wait for clk_period;
        A <= "10100110";
        B <= "01001010";
        C <= "00111010";
        wait for clk_period;
        A <= "00111101";
        B <= "10011100";
        C <= "01011000";
        wait for clk_period;
        A <= "01001101";
        B <= "01011101";
        C <= "11010010";
        wait for clk_period;
        A <= "11111011";
        B <= "10010101";
        C <= "11001111";
        wait for clk_period;
        A <= "01010001";
        B <= "00001100";
        C <= "11101101";
        wait for clk_period;
        A <= "10100111";
        B <= "10100011";
        C <= "01010001";
        wait for clk_period;
        A <= "01100001";
        B <= "01000001";
        C <= "10000111";
        wait for clk_period;
        A <= "01000101";
        B <= "01111000";
        C <= "11000111";
        wait for clk_period;
        A <= "01010000";
        B <= "01100011";
        C <= "10111110";
        wait for clk_period;
        A <= "00010010";
        B <= "11100110";
        C <= "01011111";
        wait for clk_period;
        A <= "01010001";
        B <= "10001101";
        C <= "11001011";
        wait for clk_period;
        A <= "11011100";
        B <= "01101000";
        C <= "10010111";
        wait for clk_period;
        A <= "10011110";
        B <= "10101111";
        C <= "01001001";
        wait for clk_period;
        A <= "11110110";
        B <= "01011000";
        C <= "10111001";
        wait for clk_period;
        A <= "00001100";
        B <= "11101111";
        C <= "00000111";
        wait for clk_period;
        A <= "11100101";
        B <= "01110001";
        C <= "01110111";
        wait for clk_period;
        A <= "10101110";
        B <= "01110100";
        C <= "01101101";
        wait for clk_period;
        A <= "10110110";
        B <= "10001011";
        C <= "01111110";
        wait for clk_period;
        A <= "11001110";
        B <= "11100111";
        C <= "10010100";
        wait for clk_period;
        A <= "11001000";
        B <= "11100110";
        C <= "01000101";
        wait for clk_period;
        A <= "11000111";
        B <= "00111100";
        C <= "00101011";
        wait for clk_period;
        A <= "00101000";
        B <= "01001001";
        C <= "10010111";
        wait for clk_period;
        A <= "10100010";
        B <= "11001101";
        C <= "11010000";
        wait for clk_period;
        A <= "10001100";
        B <= "00000000";
        C <= "00000110";
        wait for clk_period;
        A <= "10001101";
        B <= "10010100";
        C <= "11111011";
        wait for clk_period;
        A <= "00111101";
        B <= "01100100";
        C <= "01000010";
        wait for clk_period;
        A <= "00100100";
        B <= "10000111";
        C <= "00000001";
        wait for clk_period;
        A <= "11101110";
        B <= "00101111";
        C <= "00110110";
        wait for clk_period;
        A <= "11001100";
        B <= "01100011";
        C <= "11111100";
        wait for clk_period;
        A <= "01110000";
        B <= "00111111";
        C <= "11110110";
        wait for clk_period;
        A <= "00010110";
        B <= "11111000";
        C <= "00010100";
        wait for clk_period;
        A <= "00101110";
        B <= "10111110";
        C <= "01011100";
        wait for clk_period;
        A <= "00001001";
        B <= "11011100";
        C <= "11101011";
        wait for clk_period;
        A <= "01100111";
        B <= "00010011";
        C <= "11001100";
        wait for clk_period;
        A <= "00010110";
        B <= "00011111";
        C <= "01010000";
        wait for clk_period;
        A <= "01101011";
        B <= "11001011";
        C <= "01001000";
        wait for clk_period;
        A <= "01111110";
        B <= "00100000";
        C <= "00100000";
        wait for clk_period;
        A <= "01010100";
        B <= "01001111";
        C <= "10110010";
        wait for clk_period;
        A <= "01001000";
        B <= "10000001";
        C <= "10011010";
        wait for clk_period;
        A <= "01000111";
        B <= "00110111";
        C <= "11110001";
        wait for clk_period;
        A <= "00000110";
        B <= "00110101";
        C <= "00110101";
        wait for clk_period;
        A <= "11000110";
        B <= "11111111";
        C <= "00001011";
        wait for clk_period;
        A <= "01011101";
        B <= "00110000";
        C <= "00100111";
        wait for clk_period;
        A <= "00111111";
        B <= "00100001";
        C <= "11100010";
        wait for clk_period;
        A <= "00110100";
        B <= "00111101";
        C <= "00001001";
        wait for clk_period;
        A <= "00110011";
        B <= "00011111";
        C <= "01101011";
        wait for clk_period;
        A <= "10100000";
        B <= "10000101";
        C <= "01011100";
        wait for clk_period;
        A <= "01100000";
        B <= "01100010";
        C <= "11110000";
        wait for clk_period;
        A <= "10101100";
        B <= "11111010";
        C <= "00111101";
        wait for clk_period;
        A <= "01011110";
        B <= "11111110";
        C <= "11100101";
        wait for clk_period;
        A <= "11111100";
        B <= "10010011";
        C <= "00001010";
        wait for clk_period;
        A <= "10111100";
        B <= "01100010";
        C <= "11001100";
        wait for clk_period;
        A <= "01100001";
        B <= "00111100";
        C <= "11100110";
        wait for clk_period;
        A <= "10101001";
        B <= "10101010";
        C <= "10000001";
        wait for clk_period;
        A <= "00001001";
        B <= "11001000";
        C <= "10100010";
        wait for clk_period;
        A <= "10100001";
        B <= "11001111";
        C <= "01010001";
        wait for clk_period;
        A <= "10111011";
        B <= "10111111";
        C <= "01000100";
        wait for clk_period;
        A <= "10101001";
        B <= "10000110";
        C <= "10000000";
        wait for clk_period;
        A <= "10000011";
        B <= "01011100";
        C <= "00110000";
        wait for clk_period;
        A <= "00101001";
        B <= "01011000";
        C <= "11101100";
        wait for clk_period;
        A <= "01010010";
        B <= "00011011";
        C <= "00101100";
        wait for clk_period;
        A <= "01001010";
        B <= "11101011";
        C <= "10111001";
        wait for clk_period;
        A <= "01111001";
        B <= "00001011";
        C <= "10101011";
        wait for clk_period;
        A <= "00111111";
        B <= "10111101";
        C <= "11001011";
        wait for clk_period;
        A <= "11100101";
        B <= "11111011";
        C <= "11110001";
        wait for clk_period;
        A <= "00001111";
        B <= "11011101";
        C <= "01101101";
        wait for clk_period;
        A <= "10101110";
        B <= "01101100";
        C <= "11101001";
        wait for clk_period;
        A <= "01000001";
        B <= "11010101";
        C <= "00001110";
        wait for clk_period;
        A <= "00000110";
        B <= "01000101";
        C <= "01001111";
        wait for clk_period;
        A <= "10011000";
        B <= "11011001";
        C <= "10010010";
        wait for clk_period;
        A <= "11110011";
        B <= "01010100";
        C <= "11110110";
        wait for clk_period;
        A <= "11001000";
        B <= "11101000";
        C <= "01110011";
        wait for clk_period;
        A <= "10001011";
        B <= "11010100";
        C <= "01011000";
        wait for clk_period;
        A <= "01101101";
        B <= "01101100";
        C <= "10100000";
        wait for clk_period;
        A <= "00000110";
        B <= "10111010";
        C <= "10110110";
        wait for clk_period;
        A <= "10000000";
        B <= "01101110";
        C <= "01100001";
        wait for clk_period;
        A <= "11101111";
        B <= "01110100";
        C <= "01011101";
        wait for clk_period;
        A <= "11101111";
        B <= "00101011";
        C <= "01100000";
        wait for clk_period;
        A <= "10100100";
        B <= "01011100";
        C <= "11101100";
        wait for clk_period;
        A <= "01001001";
        B <= "10100010";
        C <= "01001010";
        wait for clk_period;
        A <= "11000110";
        B <= "00101000";
        C <= "10011100";
        wait for clk_period;
        A <= "01101010";
        B <= "10000101";
        C <= "00010010";
        wait for clk_period;
        A <= "01111001";
        B <= "00010001";
        C <= "01001101";
        wait for clk_period;
        A <= "11101110";
        B <= "00011101";
        C <= "01100111";
        wait for clk_period;
        A <= "01101011";
        B <= "10100000";
        C <= "11101000";
        wait for clk_period;
        A <= "01010110";
        B <= "00010111";
        C <= "10110000";
        wait for clk_period;
        A <= "11010100";
        B <= "11111010";
        C <= "01100001";
        wait for clk_period;
        A <= "00110111";
        B <= "00110011";
        C <= "11101011";
        wait for clk_period;
        A <= "10100010";
        B <= "00001101";
        C <= "10111010";
        wait for clk_period;
        A <= "01000011";
        B <= "01111011";
        C <= "01011101";
        wait for clk_period;
        A <= "10111001";
        B <= "11101010";
        C <= "00001111";
        wait for clk_period;
        A <= "11001001";
        B <= "11101010";
        C <= "10100111";
        wait for clk_period;
        A <= "11111100";
        B <= "11110111";
        C <= "01111011";
        wait for clk_period;
        A <= "11111011";
        B <= "00001110";
        C <= "11111101";
        wait for clk_period;
        A <= "01011010";
        B <= "00011111";
        C <= "00110001";
        wait for clk_period;
        A <= "01010110";
        B <= "10000000";
        C <= "11100000";
        wait for clk_period;
        A <= "10100010";
        B <= "01110110";
        C <= "11110010";
        wait for clk_period;
        A <= "00111111";
        B <= "11101110";
        C <= "01011000";
        wait for clk_period;
        A <= "10000011";
        B <= "00110111";
        C <= "01101000";
        wait for clk_period;
        A <= "01000101";
        B <= "01100010";
        C <= "11111100";
        wait for clk_period;
        A <= "00001000";
        B <= "11110101";
        C <= "00101100";
        wait for clk_period;
        A <= "00001101";
        B <= "00110010";
        C <= "01011110";
        wait for clk_period;
        A <= "00111011";
        B <= "01000000";
        C <= "10100110";
        wait for clk_period;
        A <= "01110001";
        B <= "10111100";
        C <= "00011110";
        wait for clk_period;
        A <= "11011011";
        B <= "01010000";
        C <= "00000111";
        wait for clk_period;
        A <= "00000001";
        B <= "00010000";
        C <= "11001101";
        wait for clk_period;
        A <= "01001100";
        B <= "10000101";
        C <= "00001110";
        wait for clk_period;
        A <= "01101101";
        B <= "10101010";
        C <= "11011000";
        wait for clk_period;
        A <= "01010011";
        B <= "00111100";
        C <= "10000110";
        wait for clk_period;
        A <= "01110011";
        B <= "10111010";
        C <= "11100001";
        wait for clk_period;
        A <= "00011010";
        B <= "01000010";
        C <= "11100111";
        wait for clk_period;
        A <= "00010111";
        B <= "11111001";
        C <= "01110100";
        wait for clk_period;
        A <= "10110010";
        B <= "10001000";
        C <= "11111101";
        wait for clk_period;
        A <= "10100000";
        B <= "11111111";
        C <= "00100101";
        wait for clk_period;
        A <= "01011110";
        B <= "11111101";
        C <= "01101100";
        wait for clk_period;
        A <= "01101000";
        B <= "11110100";
        C <= "11101010";
        wait for clk_period;
        A <= "00000001";
        B <= "01011110";
        C <= "10001000";
        wait for clk_period;
        A <= "10001011";
        B <= "00001111";
        C <= "00100111";
        wait for clk_period;
        A <= "11001100";
        B <= "10101000";
        C <= "10001000";
        wait for clk_period;
        A <= "10000000";
        B <= "11110010";
        C <= "01110110";
        wait for clk_period;
        A <= "10100100";
        B <= "11110111";
        C <= "10111100";
        wait for clk_period;
        A <= "01001000";
        B <= "10111110";
        C <= "01010010";
        wait for clk_period;
        A <= "11011111";
        B <= "00110000";
        C <= "11110011";
        wait for clk_period;
        A <= "00111100";
        B <= "10011001";
        C <= "00100110";
        wait for clk_period;
        A <= "11001100";
        B <= "01011101";
        C <= "00100101";
        wait for clk_period;
        A <= "10101001";
        B <= "11010101";
        C <= "00100011";
        wait for clk_period;
        A <= "11101000";
        B <= "00000011";
        C <= "11111100";
        wait for clk_period;
        A <= "00010010";
        B <= "00100011";
        C <= "00001011";
        wait for clk_period;
        A <= "00111011";
        B <= "00100101";
        C <= "01100011";
        wait for clk_period;
        A <= "11001100";
        B <= "10011101";
        C <= "00010110";
        wait for clk_period;
        A <= "01100011";
        B <= "01010110";
        C <= "00101000";
        wait for clk_period;
        A <= "01101010";
        B <= "00101110";
        C <= "10010101";
        wait for clk_period;
        A <= "10111000";
        B <= "01011110";
        C <= "10001111";
        wait for clk_period;
        A <= "10110101";
        B <= "01100001";
        C <= "10010010";
        wait for clk_period;
        A <= "11101110";
        B <= "10001000";
        C <= "00111100";
        wait for clk_period;
        A <= "00100000";
        B <= "11010011";
        C <= "00111110";
        wait for clk_period;
        A <= "00001001";
        B <= "01110010";
        C <= "01111100";
        wait for clk_period;
        A <= "00011100";
        B <= "00010011";
        C <= "11000000";
        wait for clk_period;
        A <= "11111000";
        B <= "10010110";
        C <= "01100000";
        wait for clk_period;
        A <= "01100011";
        B <= "10011010";
        C <= "10001001";
        wait for clk_period;
        A <= "10011010";
        B <= "10100111";
        C <= "11011100";
        wait for clk_period;
        A <= "01111001";
        B <= "01101010";
        C <= "11011011";
        wait for clk_period;
        A <= "10010011";
        B <= "01011110";
        C <= "11011010";
        wait for clk_period;
        A <= "10001111";
        B <= "11010001";
        C <= "00010000";
        wait for clk_period;
        A <= "01110111";
        B <= "01101011";
        C <= "01000001";
        wait for clk_period;
        A <= "01000011";
        B <= "10100111";
        C <= "10100100";
        wait for clk_period;
        A <= "10010011";
        B <= "01001000";
        C <= "00110101";
        wait for clk_period;
        A <= "00000010";
        B <= "01010010";
        C <= "01011110";
        wait for clk_period;
        A <= "11010100";
        B <= "00010011";
        C <= "10111101";
        wait for clk_period;
        A <= "01110111";
        B <= "01010100";
        C <= "11101101";
        wait for clk_period;
        A <= "10110111";
        B <= "10001110";
        C <= "01000010";
        wait for clk_period;
        A <= "00000011";
        B <= "10011010";
        C <= "00111000";
        wait for clk_period;
        A <= "11000111";
        B <= "01011100";
        C <= "11010010";
        wait for clk_period;
        A <= "11101100";
        B <= "01010011";
        C <= "01010110";
        wait for clk_period;
        A <= "01110100";
        B <= "00000011";
        C <= "11100111";
        wait for clk_period;
        A <= "10010101";
        B <= "00001111";
        C <= "11010110";
        wait for clk_period;
        A <= "10010011";
        B <= "10000000";
        C <= "01001101";
        wait for clk_period;
        A <= "00101101";
        B <= "10011011";
        C <= "11010011";
        wait for clk_period;
        A <= "01010010";
        B <= "11001100";
        C <= "00101010";
        wait for clk_period;
        A <= "00001001";
        B <= "11000100";
        C <= "10011111";
        wait for clk_period;
        A <= "00111000";
        B <= "01000011";
        C <= "11000110";
        wait for clk_period;
        A <= "01101111";
        B <= "00100111";
        C <= "00000110";
        wait for clk_period;
        A <= "01011110";
        B <= "11011001";
        C <= "11010110";
        wait for clk_period;
        A <= "10001101";
        B <= "11011101";
        C <= "10111110";
        wait for clk_period;
        A <= "11010111";
        B <= "11111110";
        C <= "11110010";
        wait for clk_period;
        A <= "00111011";
        B <= "11110011";
        C <= "00001001";
        wait for clk_period;
        A <= "01100111";
        B <= "11110100";
        C <= "10011100";
        wait for clk_period;
        A <= "00111001";
        B <= "10000110";
        C <= "11000111";
        wait for clk_period;
        A <= "01010111";
        B <= "11011010";
        C <= "10101001";
        wait for clk_period;
        A <= "01000110";
        B <= "00011001";
        C <= "10010000";
        wait for clk_period;
        A <= "10110000";
        B <= "01110010";
        C <= "01011100";
        wait for clk_period;
        A <= "11000000";
        B <= "00000011";
        C <= "00000100";
        wait for clk_period;
        A <= "11001110";
        B <= "01000110";
        C <= "10011011";
        wait for clk_period;
        A <= "01010111";
        B <= "00011101";
        C <= "00101100";
        wait for clk_period;
        A <= "00100111";
        B <= "01111110";
        C <= "00010111";
        wait for clk_period;
        A <= "10001100";
        B <= "11101010";
        C <= "10010100";
        wait for clk_period;
        A <= "10110000";
        B <= "01111111";
        C <= "11011111";
        wait for clk_period;
        A <= "00110101";
        B <= "11011111";
        C <= "10000101";
        wait for clk_period;
        A <= "10111010";
        B <= "01001011";
        C <= "01011111";
        wait for clk_period;
        A <= "01110101";
        B <= "01101101";
        C <= "10010101";
        wait for clk_period;
        A <= "01110011";
        B <= "01100110";
        C <= "11100110";
        wait for clk_period;
        A <= "10100010";
        B <= "01000001";
        C <= "01111111";
        wait for clk_period;
        A <= "01111011";
        B <= "01110011";
        C <= "11111101";
        wait for clk_period;
        A <= "00110110";
        B <= "00100001";
        C <= "11110111";
        wait for clk_period;
        A <= "01101111";
        B <= "11101110";
        C <= "01010001";
        wait for clk_period;
        A <= "11000000";
        B <= "01100100";
        C <= "01000111";
        wait for clk_period;
        A <= "01010101";
        B <= "10011111";
        C <= "01011101";
        wait for clk_period;
        A <= "11111011";
        B <= "10100111";
        C <= "00111000";
        wait for clk_period;
        A <= "00010111";
        B <= "00010011";
        C <= "11101011";
        wait for clk_period;
        A <= "10011101";
        B <= "01011001";
        C <= "00001111";
        wait for clk_period;
        A <= "00110110";
        B <= "00110000";
        C <= "01110011";
        wait for clk_period;
        A <= "11111100";
        B <= "10111000";
        C <= "11000010";
        wait for clk_period;
        A <= "11111010";
        B <= "00101101";
        C <= "01000101";
        wait for clk_period;
        A <= "01110001";
        B <= "10010110";
        C <= "00111011";
        wait for clk_period;
        A <= "01010000";
        B <= "10101100";
        C <= "00110000";
        wait for clk_period;
        A <= "11001011";
        B <= "00100100";
        C <= "00111011";
        wait for clk_period;
        A <= "10000101";
        B <= "01111110";
        C <= "01111000";
        wait for clk_period;
        A <= "01100111";
        B <= "11101100";
        C <= "01100111";
        wait for clk_period;
        A <= "10111101";
        B <= "01011100";
        C <= "11111000";
        wait for clk_period;
        A <= "11001110";
        B <= "10110011";
        C <= "00110001";
        wait for clk_period;
        A <= "11110011";
        B <= "10101000";
        C <= "11111101";
        wait for clk_period;
        A <= "00110001";
        B <= "00000010";
        C <= "01010011";
        wait for clk_period;
        A <= "11011111";
        B <= "01110001";
        C <= "01101111";
        wait for clk_period;
        A <= "01111010";
        B <= "10110100";
        C <= "01001101";
        wait for clk_period;
        A <= "01010101";
        B <= "11101011";
        C <= "00111101";
        wait for clk_period;
        A <= "01111010";
        B <= "10000110";
        C <= "10011101";
        wait for clk_period;
        A <= "00101111";
        B <= "00111001";
        C <= "11111000";
        wait for clk_period;
        A <= "00000100";
        B <= "11011011";
        C <= "01111000";
        wait for clk_period;
        A <= "10000000";
        B <= "10100101";
        C <= "11010111";
        wait for clk_period;
        A <= "10010010";
        B <= "00110010";
        C <= "00111101";
        wait for clk_period;
        A <= "01111010";
        B <= "01011111";
        C <= "10101000";
        wait for clk_period;
        A <= "11010001";
        B <= "00111101";
        C <= "01000000";
        wait for clk_period;
        A <= "00011101";
        B <= "11101011";
        C <= "01111000";
        wait for clk_period;
        A <= "10010001";
        B <= "01110010";
        C <= "01001101";
        wait for clk_period;
        A <= "10011100";
        B <= "10111011";
        C <= "00111110";
        wait for clk_period;
        A <= "10000000";
        B <= "00100011";
        C <= "00000101";
        wait for clk_period;
        A <= "10000000";
        B <= "10110000";
        C <= "11001110";
        wait for clk_period;
        A <= "11110101";
        B <= "11110110";
        C <= "10001000";
        wait for clk_period;
        A <= "00011011";
        B <= "10111000";
        C <= "11100010";
        wait for clk_period;
        A <= "01101001";
        B <= "11011111";
        C <= "01011110";
        wait for clk_period;
        A <= "11110011";
        B <= "10111010";
        C <= "11101011";
        wait for clk_period;
        A <= "10001001";
        B <= "10010000";
        C <= "00001011";
        wait for clk_period;
        A <= "01100010";
        B <= "11110010";
        C <= "11111101";
        wait for clk_period;
        A <= "00000001";
        B <= "10001101";
        C <= "00100110";
        wait for clk_period;
        A <= "11000000";
        B <= "11111000";
        C <= "00011001";
        wait for clk_period;
        A <= "11000001";
        B <= "11001001";
        C <= "01101101";
        wait for clk_period;
        A <= "11010110";
        B <= "01000100";
        C <= "00001011";
        wait for clk_period;
        A <= "01010010";
        B <= "10000011";
        C <= "01010001";
        wait for clk_period;
        A <= "10101011";
        B <= "10011000";
        C <= "01001101";
        wait for clk_period;
        A <= "00101110";
        B <= "00110100";
        C <= "11110110";
        wait for clk_period;
        A <= "11011000";
        B <= "11011011";
        C <= "10011010";
        wait for clk_period;
        A <= "10000011";
        B <= "01000100";
        C <= "10110100";
        wait for clk_period;
        A <= "00011001";
        B <= "01000101";
        C <= "11000101";
        wait for clk_period;
        A <= "11011001";
        B <= "10011110";
        C <= "10100000";
        wait for clk_period;
        A <= "11100111";
        B <= "11001111";
        C <= "01110100";
        wait for clk_period;
        A <= "00010011";
        B <= "10011100";
        C <= "00010001";
        wait for clk_period;
        A <= "01100000";
        B <= "11110011";
        C <= "11000101";
        wait for clk_period;
        A <= "10100111";
        B <= "10010100";
        C <= "10001111";
        wait for clk_period;
        A <= "10111010";
        B <= "11000010";
        C <= "01111010";
        wait for clk_period;
        A <= "00000111";
        B <= "11000100";
        C <= "10001111";
        wait for clk_period;
        A <= "11110010";
        B <= "00100100";
        C <= "10010100";
        wait for clk_period;
        A <= "10110011";
        B <= "11011011";
        C <= "01100100";
        wait for clk_period;
        A <= "10001111";
        B <= "00011001";
        C <= "10000000";
        wait for clk_period;
        A <= "10101010";
        B <= "11001011";
        C <= "11110100";
        wait for clk_period;
        A <= "00111010";
        B <= "01111000";
        C <= "10100010";
        wait for clk_period;
        A <= "00100110";
        B <= "10000011";
        C <= "01001011";
        wait for clk_period;
        A <= "00110010";
        B <= "10100100";
        C <= "00111010";
        wait for clk_period;
        A <= "11000001";
        B <= "10010010";
        C <= "10100100";
        wait for clk_period;
        A <= "00110010";
        B <= "10111110";
        C <= "01100000";
        wait for clk_period;
        A <= "01001110";
        B <= "11000100";
        C <= "10001001";
        wait for clk_period;
        A <= "00110000";
        B <= "00011100";
        C <= "10001111";
        wait for clk_period;
        A <= "01000010";
        B <= "11010111";
        C <= "10001001";
        wait for clk_period;
        A <= "01110011";
        B <= "00001000";
        C <= "11110001";
        wait for clk_period;
        A <= "00001010";
        B <= "00001010";
        C <= "10111001";
        wait for clk_period;
        A <= "00111111";
        B <= "00101111";
        C <= "11011000";
        wait for clk_period;
        A <= "11010101";
        B <= "01010111";
        C <= "11101011";
        wait for clk_period;
        A <= "10011001";
        B <= "11110111";
        C <= "10011011";
        wait for clk_period;
        A <= "00001100";
        B <= "00001001";
        C <= "01111011";
        wait for clk_period;
        A <= "00101000";
        B <= "10100110";
        C <= "00001000";
        wait for clk_period;
        A <= "01111010";
        B <= "10000001";
        C <= "11011100";
        wait for clk_period;
        A <= "10101001";
        B <= "00000111";
        C <= "11010111";
        wait for clk_period;
        A <= "01011101";
        B <= "00111000";
        C <= "11001111";
        wait for clk_period;
        A <= "01100011";
        B <= "00010001";
        C <= "10110001";
        wait for clk_period;
        A <= "00111001";
        B <= "10101101";
        C <= "11000010";
        wait for clk_period;
        A <= "11110100";
        B <= "01001111";
        C <= "01001000";
        wait for clk_period;
        A <= "11011000";
        B <= "11010001";
        C <= "11100011";
        wait for clk_period;
        A <= "00010011";
        B <= "11110100";
        C <= "00111110";
        wait for clk_period;
        A <= "10101000";
        B <= "00001111";
        C <= "01100111";
        wait for clk_period;
        A <= "01111000";
        B <= "11110000";
        C <= "01001001";
        wait for clk_period;
        A <= "11000100";
        B <= "01110000";
        C <= "01110111";
        wait for clk_period;
        A <= "00100011";
        B <= "01000101";
        C <= "10100101";
        wait for clk_period;
        A <= "11000101";
        B <= "00111001";
        C <= "10100000";
        wait for clk_period;
        A <= "01111010";
        B <= "00011010";
        C <= "10011100";
        wait for clk_period;
        A <= "10100000";
        B <= "11011011";
        C <= "11000011";
        wait for clk_period;
        A <= "01001000";
        B <= "10010100";
        C <= "00101001";
        wait for clk_period;
        A <= "10101001";
        B <= "11011110";
        C <= "10011110";
        wait for clk_period;
        A <= "00100001";
        B <= "10111011";
        C <= "01100111";
        wait for clk_period;
        A <= "00110010";
        B <= "00100100";
        C <= "10000001";
        wait for clk_period;
        A <= "00111111";
        B <= "10111011";
        C <= "01001111";
        wait for clk_period;
        A <= "10010100";
        B <= "01000110";
        C <= "11001100";
        wait for clk_period;
        A <= "10111011";
        B <= "01001100";
        C <= "01110010";
        wait for clk_period;
        A <= "11110010";
        B <= "01010111";
        C <= "11001011";
        wait for clk_period;
        A <= "01111111";
        B <= "11011101";
        C <= "10111010";
        wait for clk_period;
        A <= "00011011";
        B <= "01011101";
        C <= "00111011";
        wait for clk_period;
        A <= "00110110";
        B <= "01100101";
        C <= "11011111";
        wait for clk_period;
        A <= "00110010";
        B <= "01000101";
        C <= "11001001";
        wait for clk_period;
        A <= "11101011";
        B <= "00010100";
        C <= "01000101";
        wait for clk_period;
        A <= "00101000";
        B <= "01010110";
        C <= "11100111";
        wait for clk_period;
        A <= "00001001";
        B <= "11110001";
        C <= "00111101";
        wait for clk_period;
        A <= "00000100";
        B <= "10100101";
        C <= "01111100";
        wait for clk_period;
        A <= "11110100";
        B <= "10000100";
        C <= "10010101";
        wait for clk_period;
        A <= "11011100";
        B <= "10111001";
        C <= "11101100";
        wait for clk_period;
        A <= "01111111";
        B <= "11110111";
        C <= "00110001";
        wait for clk_period;
        A <= "00011100";
        B <= "01000101";
        C <= "00111000";
        wait for clk_period;
        A <= "11100100";
        B <= "00110110";
        C <= "00001000";
        wait for clk_period;
        A <= "10010110";
        B <= "01000100";
        C <= "01011110";
        wait for clk_period;
        A <= "10001101";
        B <= "10101110";
        C <= "11001011";
        wait for clk_period;
        A <= "00001101";
        B <= "10000010";
        C <= "01110010";
        wait for clk_period;
        A <= "01010001";
        B <= "10001110";
        C <= "01000111";
        wait for clk_period;
        A <= "10011101";
        B <= "11110100";
        C <= "11100101";
        wait for clk_period;
        A <= "10010011";
        B <= "11101110";
        C <= "01011100";
        wait for clk_period;
        A <= "11010110";
        B <= "00101011";
        C <= "00111111";
        wait for clk_period;
        A <= "00100100";
        B <= "00110111";
        C <= "10101100";
        wait for clk_period;
        A <= "00111000";
        B <= "11101010";
        C <= "00011101";
        wait for clk_period;
        A <= "01100111";
        B <= "00101000";
        C <= "10010011";
        wait for clk_period;
        A <= "11000111";
        B <= "00111011";
        C <= "00010111";
        wait for clk_period;
        A <= "01100111";
        B <= "00101011";
        C <= "00111001";
        wait for clk_period;
        A <= "00100101";
        B <= "11011100";
        C <= "01001001";
        wait for clk_period;
        A <= "00110011";
        B <= "01000101";
        C <= "11100010";
        wait for clk_period;
        A <= "10110111";
        B <= "01111000";
        C <= "10001001";
        wait for clk_period;
        A <= "11111101";
        B <= "10010011";
        C <= "11011000";
        wait for clk_period;
        A <= "11001000";
        B <= "01110010";
        C <= "11000100";
        wait for clk_period;
        A <= "01000101";
        B <= "11100011";
        C <= "00001010";
        wait for clk_period;
        A <= "10111100";
        B <= "01010001";
        C <= "00111111";
        wait for clk_period;
        A <= "11110000";
        B <= "11101110";
        C <= "10000011";
        wait for clk_period;
        A <= "10110011";
        B <= "01100001";
        C <= "01101101";
        wait for clk_period;
        A <= "11110000";
        B <= "11010011";
        C <= "01100111";
        wait for clk_period;
        A <= "11111000";
        B <= "01100111";
        C <= "10100110";
        wait for clk_period;
        A <= "00010110";
        B <= "11001000";
        C <= "10010110";
        wait for clk_period;
        A <= "11010011";
        B <= "10010100";
        C <= "11100100";
        wait for clk_period;
        A <= "10101101";
        B <= "11010101";
        C <= "00110101";
        wait for clk_period;
        A <= "10101101";
        B <= "01011000";
        C <= "10010001";
        wait for clk_period;
        A <= "00100111";
        B <= "01001101";
        C <= "00000101";
        wait for clk_period;
        A <= "00001111";
        B <= "11110100";
        C <= "00010101";
        wait for clk_period;
        A <= "10000110";
        B <= "11010010";
        C <= "00101001";
        wait for clk_period;
        A <= "11100011";
        B <= "01001100";
        C <= "10111011";
        wait for clk_period;
        A <= "00110000";
        B <= "00100001";
        C <= "01101010";
        wait for clk_period;
        A <= "10111010";
        B <= "01000100";
        C <= "00001010";
        wait for clk_period;
        A <= "00101111";
        B <= "00011000";
        C <= "00111010";
        wait for clk_period;
        A <= "11110010";
        B <= "00011000";
        C <= "01101001";
        wait for clk_period;
        A <= "01110011";
        B <= "00110000";
        C <= "11110111";
        wait for clk_period;
        A <= "01011110";
        B <= "01001011";
        C <= "11011000";
        wait for clk_period;
        A <= "10010000";
        B <= "10110100";
        C <= "01101111";
        wait for clk_period;
        A <= "01100110";
        B <= "00100001";
        C <= "11111100";
        wait for clk_period;
        A <= "01000100";
        B <= "10111011";
        C <= "00101010";
        wait for clk_period;
        A <= "11011001";
        B <= "01101010";
        C <= "00110001";
        wait for clk_period;
        A <= "00001100";
        B <= "01101010";
        C <= "10111011";
        wait for clk_period;
        A <= "00000110";
        B <= "11000010";
        C <= "11011010";
        wait for clk_period;
        A <= "11111101";
        B <= "00000010";
        C <= "11011110";
        wait for clk_period;
        A <= "00000001";
        B <= "01110010";
        C <= "10001110";
        wait for clk_period;
        A <= "01101011";
        B <= "11011011";
        C <= "01100100";
        wait for clk_period;
        A <= "11100101";
        B <= "10110100";
        C <= "11001001";
        wait for clk_period;
        A <= "00101110";
        B <= "11000110";
        C <= "00010110";
        wait for clk_period;
        A <= "10100110";
        B <= "00000011";
        C <= "10110111";
        wait for clk_period;
        A <= "10111101";
        B <= "00101111";
        C <= "00010101";
        wait for clk_period;
        A <= "11011010";
        B <= "11111010";
        C <= "11011010";
        wait for clk_period;
        A <= "11110001";
        B <= "01001010";
        C <= "01111000";
        wait for clk_period;
        A <= "11010100";
        B <= "00111110";
        C <= "11101111";
        wait for clk_period;
        A <= "11111111";
        B <= "01001110";
        C <= "01010011";
        wait for clk_period;
        A <= "11111100";
        B <= "10010000";
        C <= "10110000";
        wait for clk_period;
        A <= "11100010";
        B <= "01001000";
        C <= "01011000";
        wait for clk_period;
        A <= "00110110";
        B <= "10000101";
        C <= "00101011";
        wait for clk_period;
        A <= "01000110";
        B <= "10010000";
        C <= "10111001";
        wait for clk_period;
        A <= "11011000";
        B <= "00001010";
        C <= "00100101";
        wait for clk_period;
        A <= "00100110";
        B <= "00010000";
        C <= "01010110";
        wait for clk_period;
        A <= "10110011";
        B <= "10101100";
        C <= "01101100";
        wait for clk_period;
        A <= "01101101";
        B <= "10101110";
        C <= "10100001";
        wait for clk_period;
        A <= "11101100";
        B <= "11011111";
        C <= "00000100";
        wait for clk_period;
        A <= "00011110";
        B <= "11011101";
        C <= "01101101";
        wait for clk_period;
        A <= "01010110";
        B <= "10111100";
        C <= "00011001";
        wait for clk_period;
        A <= "00111000";
        B <= "10001011";
        C <= "01001110";
        wait for clk_period;
        A <= "11111000";
        B <= "01100101";
        C <= "01100100";
        wait for clk_period;
        A <= "10100101";
        B <= "00010110";
        C <= "10111001";
        wait for clk_period;
        A <= "11110110";
        B <= "00111101";
        C <= "00001100";
        wait for clk_period;
        A <= "00001110";
        B <= "00011101";
        C <= "00011110";
        wait for clk_period;
        A <= "11111101";
        B <= "01001111";
        C <= "00100011";
        wait for clk_period;
        A <= "11101001";
        B <= "01010111";
        C <= "11000000";
        wait for clk_period;
        A <= "10111010";
        B <= "10110100";
        C <= "10000111";
        wait for clk_period;
        A <= "10111100";
        B <= "01010011";
        C <= "10100101";
        wait for clk_period;
        A <= "01011011";
        B <= "11011010";
        C <= "01101111";
        wait for clk_period;
        A <= "11000000";
        B <= "01111110";
        C <= "00100110";
        wait for clk_period;
        A <= "01001110";
        B <= "10110111";
        C <= "01011000";
        wait for clk_period;
        A <= "10111111";
        B <= "00000011";
        C <= "11111101";
        wait for clk_period;
        A <= "10011100";
        B <= "00111010";
        C <= "11111010";
        wait for clk_period;
        A <= "00101011";
        B <= "01001000";
        C <= "11010001";
        wait for clk_period;
        A <= "01001100";
        B <= "10000010";
        C <= "10011000";
        wait for clk_period;
        A <= "00100110";
        B <= "11111010";
        C <= "10010000";
        wait for clk_period;
        A <= "10101100";
        B <= "10001001";
        C <= "01010011";
        wait for clk_period;
        A <= "10001111";
        B <= "01000110";
        C <= "10111010";
        wait for clk_period;
        A <= "01100001";
        B <= "10001000";
        C <= "11100001";
        wait for clk_period;
        A <= "00001001";
        B <= "11011010";
        C <= "11011011";
        wait for clk_period;
        A <= "01110100";
        B <= "00101011";
        C <= "00100100";
        wait for clk_period;
        A <= "10000110";
        B <= "11000010";
        C <= "00011111";
        wait for clk_period;
        A <= "00000100";
        B <= "00000111";
        C <= "10110000";
        wait for clk_period;
        A <= "11111111";
        B <= "01101010";
        C <= "10100101";
        wait for clk_period;
        A <= "00100110";
        B <= "10101100";
        C <= "01100010";
        wait for clk_period;
        A <= "11101100";
        B <= "11010100";
        C <= "00100101";
        wait for clk_period;
        A <= "01110111";
        B <= "11111010";
        C <= "00111000";
        wait for clk_period;
        A <= "10100101";
        B <= "01101011";
        C <= "10011001";
        wait for clk_period;
        A <= "10111010";
        B <= "00001100";
        C <= "00001000";
        wait for clk_period;
        A <= "11010011";
        B <= "01000000";
        C <= "01101011";
        wait for clk_period;
        A <= "10111110";
        B <= "11111001";
        C <= "01111011";
        wait for clk_period;
        A <= "10011000";
        B <= "01101101";
        C <= "01001010";
        wait for clk_period;
        A <= "10011011";
        B <= "00011101";
        C <= "11000010";
        wait for clk_period;
        A <= "11101001";
        B <= "10010001";
        C <= "01010010";
        wait for clk_period;
        A <= "11001100";
        B <= "00110101";
        C <= "01111100";
        wait for clk_period;
        A <= "10100111";
        B <= "01000100";
        C <= "10010111";
        wait for clk_period;
        A <= "11100111";
        B <= "00111110";
        C <= "00010111";
        wait for clk_period;
        A <= "00011001";
        B <= "11010010";
        C <= "10101111";
        wait for clk_period;
        A <= "11110111";
        B <= "00100001";
        C <= "00101100";
        wait for clk_period;
        A <= "11011010";
        B <= "11001001";
        C <= "10001000";
        wait for clk_period;
        A <= "01101000";
        B <= "00100101";
        C <= "00111111";
        wait for clk_period;
        A <= "11101000";
        B <= "00010100";
        C <= "11010111";
        wait for clk_period;
        A <= "00100010";
        B <= "11001001";
        C <= "11011000";
        wait for clk_period;
        A <= "11111101";
        B <= "01110110";
        C <= "11011110";
        wait for clk_period;
        A <= "10111101";
        B <= "10010011";
        C <= "11010011";
        wait for clk_period;
        A <= "11100011";
        B <= "00110101";
        C <= "10111011";
        wait for clk_period;
        A <= "11011110";
        B <= "11010100";
        C <= "10011001";
        wait for clk_period;
        A <= "10101101";
        B <= "11111011";
        C <= "00001100";
        wait for clk_period;
        A <= "10011011";
        B <= "00001111";
        C <= "10100001";
        wait for clk_period;
        A <= "10000000";
        B <= "10101001";
        C <= "10101010";
        wait for clk_period;
        A <= "00001011";
        B <= "00110110";
        C <= "00111110";
        wait for clk_period;
        A <= "01100111";
        B <= "10011100";
        C <= "00100001";
        wait for clk_period;
        A <= "00011110";
        B <= "11101101";
        C <= "11111000";
        wait for clk_period;
        A <= "01101100";
        B <= "10001100";
        C <= "11110100";
        wait for clk_period;
        A <= "11000100";
        B <= "00010010";
        C <= "11011100";
        wait for clk_period;
        A <= "01010000";
        B <= "00010101";
        C <= "10101111";
        wait for clk_period;
        A <= "10011100";
        B <= "11101000";
        C <= "00001000";
        wait for clk_period;
        A <= "01111100";
        B <= "00111010";
        C <= "11111110";
        wait for clk_period;
        A <= "10100100";
        B <= "11111111";
        C <= "10001000";
        wait for clk_period;
        A <= "11100010";
        B <= "11001011";
        C <= "11100110";
        wait for clk_period;
        A <= "11001111";
        B <= "10000111";
        C <= "11001111";
        wait for clk_period;
        A <= "11011011";
        B <= "10101110";
        C <= "00001000";
        wait for clk_period;
        A <= "10011010";
        B <= "00101001";
        C <= "00110000";
        wait for clk_period;
        A <= "10011110";
        B <= "01000001";
        C <= "11001001";
        wait for clk_period;
        A <= "11010010";
        B <= "11111001";
        C <= "00111111";
        wait for clk_period;
        A <= "10011011";
        B <= "11111110";
        C <= "00011000";
        wait for clk_period;
        A <= "00011100";
        B <= "00110010";
        C <= "10001100";
        wait for clk_period;
        A <= "11010010";
        B <= "01110000";
        C <= "00000100";
        wait for clk_period;
        A <= "00000010";
        B <= "00010110";
        C <= "00110000";
        wait for clk_period;
        A <= "11101101";
        B <= "00000110";
        C <= "01100111";
        wait for clk_period;
        A <= "11110011";
        B <= "01001111";
        C <= "11000011";
        wait for clk_period;
        A <= "11010000";
        B <= "00100101";
        C <= "11000010";
        wait for clk_period;
        A <= "00111100";
        B <= "10111001";
        C <= "01101000";
        wait for clk_period;
        A <= "00000111";
        B <= "01011011";
        C <= "01010101";
        wait for clk_period;
        A <= "10010110";
        B <= "11011110";
        C <= "11111110";
        wait for clk_period;
        A <= "00000000";
        B <= "11111010";
        C <= "10100101";
        wait for clk_period;
        A <= "01101001";
        B <= "11001100";
        C <= "01111001";
        wait for clk_period;
        A <= "00100111";
        B <= "10101100";
        C <= "01111010";
        wait for clk_period;
        A <= "01101000";
        B <= "00101111";
        C <= "00110011";
        wait for clk_period;
        A <= "10010110";
        B <= "00110100";
        C <= "01011100";
        wait for clk_period;
        A <= "01000010";
        B <= "00100010";
        C <= "01000000";
        wait for clk_period;
        A <= "10100101";
        B <= "10000100";
        C <= "11101101";
        wait for clk_period;
        A <= "01101100";
        B <= "10000011";
        C <= "10011001";
        wait for clk_period;
        A <= "11000101";
        B <= "00100111";
        C <= "00001000";
        wait for clk_period;
        A <= "01000001";
        B <= "10111011";
        C <= "10101011";
        wait for clk_period;
        A <= "10110000";
        B <= "01111011";
        C <= "11000110";
        wait for clk_period;
        A <= "11011110";
        B <= "00100001";
        C <= "01001000";
        wait for clk_period;
        A <= "11100011";
        B <= "10000111";
        C <= "01100001";
        wait for clk_period;
        A <= "01100000";
        B <= "10011110";
        C <= "01110010";
        wait for clk_period;
        A <= "11010100";
        B <= "10100010";
        C <= "11010010";
        wait for clk_period;
        A <= "11010101";
        B <= "11001001";
        C <= "00101101";
        wait for clk_period;
        A <= "01011001";
        B <= "01001001";
        C <= "01011111";
        wait for clk_period;
        A <= "01001101";
        B <= "11111111";
        C <= "00011100";
        wait for clk_period;
        A <= "10101110";
        B <= "01000000";
        C <= "11000101";
        wait for clk_period;
        A <= "01111001";
        B <= "01010111";
        C <= "11110010";
        wait for clk_period;
        A <= "10111101";
        B <= "11010001";
        C <= "10011111";
        wait for clk_period;
        A <= "11101000";
        B <= "00100111";
        C <= "10101101";
        wait for clk_period;
        A <= "11100011";
        B <= "00101001";
        C <= "10101110";
        wait for clk_period;
        A <= "01101001";
        B <= "10101110";
        C <= "01100011";
        wait for clk_period;
        A <= "10110000";
        B <= "00110110";
        C <= "00111111";
        wait for clk_period;
        A <= "01111011";
        B <= "01111111";
        C <= "11111111";
        wait for clk_period;
        A <= "11100011";
        B <= "10001000";
        C <= "00011101";
        wait for clk_period;
        A <= "01111111";
        B <= "11011101";
        C <= "10011111";
        wait for clk_period;
        A <= "10000000";
        B <= "01001100";
        C <= "01110000";
        wait for clk_period;
        A <= "10000001";
        B <= "11111111";
        C <= "10001001";
        wait for clk_period;
        A <= "00000100";
        B <= "11000100";
        C <= "10010011";
        wait for clk_period;
        A <= "11110100";
        B <= "11100101";
        C <= "10010111";
        wait for clk_period;
        A <= "11001011";
        B <= "11001100";
        C <= "01011111";
        wait for clk_period;
        A <= "01010011";
        B <= "10011101";
        C <= "11111010";
        wait for clk_period;
        A <= "00111111";
        B <= "00111000";
        C <= "10010100";
        wait for clk_period;
        A <= "10110001";
        B <= "00100010";
        C <= "10000111";
        wait for clk_period;
        A <= "11100011";
        B <= "11110010";
        C <= "01110111";
        wait for clk_period;
        A <= "00001010";
        B <= "10001110";
        C <= "00111111";
        wait for clk_period;
        A <= "01110010";
        B <= "00100010";
        C <= "01001111";
        wait for clk_period;
        A <= "10110100";
        B <= "01000100";
        C <= "01100010";
        wait for clk_period;
        A <= "01011101";
        B <= "01001111";
        C <= "10100011";
        wait for clk_period;
        A <= "01101010";
        B <= "00100110";
        C <= "10101010";
        wait for clk_period;
        A <= "00011101";
        B <= "11100110";
        C <= "10000000";
        wait for clk_period;
        A <= "00011111";
        B <= "01100101";
        C <= "00010010";
        wait for clk_period;
        A <= "01100000";
        B <= "00101111";
        C <= "00010001";
        wait for clk_period;
        A <= "11010111";
        B <= "00100011";
        C <= "10100001";
        wait for clk_period;
        A <= "01111010";
        B <= "10000011";
        C <= "01100000";
        wait for clk_period;
        A <= "10100110";
        B <= "10001010";
        C <= "00100110";
        wait for clk_period;
        A <= "00111010";
        B <= "11100110";
        C <= "01101000";
        wait for clk_period;
        A <= "01011001";
        B <= "00111111";
        C <= "00010010";
        wait for clk_period;
        A <= "01100110";
        B <= "11000111";
        C <= "10011110";
        wait for clk_period;
        A <= "10110111";
        B <= "01010111";
        C <= "10110100";
        wait for clk_period;
        A <= "11110111";
        B <= "10101001";
        C <= "11001100";
        wait for clk_period;
        A <= "11101100";
        B <= "10000100";
        C <= "10101001";
        wait for clk_period;
        A <= "10010110";
        B <= "10001100";
        C <= "00000101";
        wait for clk_period;
        A <= "00000110";
        B <= "00011001";
        C <= "10101010";
        wait for clk_period;
        A <= "01011110";
        B <= "10011011";
        C <= "00100100";
        wait for clk_period;
        A <= "10110001";
        B <= "00111001";
        C <= "11110001";
        wait for clk_period;
        A <= "01100011";
        B <= "10001010";
        C <= "11111000";
        wait for clk_period;
        A <= "00110110";
        B <= "01010100";
        C <= "01001001";
        wait for clk_period;
        A <= "01000100";
        B <= "01011010";
        C <= "00001010";
        wait for clk_period;
        A <= "00001001";
        B <= "11111001";
        C <= "10100001";
        wait for clk_period;
        A <= "10011011";
        B <= "01000111";
        C <= "01011000";
        wait for clk_period;
        A <= "11001010";
        B <= "00001101";
        C <= "00111100";
        wait for clk_period;
        A <= "11111010";
        B <= "01101111";
        C <= "10100010";
        wait for clk_period;
        A <= "00110101";
        B <= "01100001";
        C <= "10000010";
        wait for clk_period;
        A <= "10010000";
        B <= "11001001";
        C <= "01001111";
        wait for clk_period;
        A <= "10001100";
        B <= "01110111";
        C <= "00101011";
        wait for clk_period;
        A <= "11010010";
        B <= "11001011";
        C <= "01111001";
        wait for clk_period;
        A <= "00010001";
        B <= "00000110";
        C <= "01100011";
        wait for clk_period;
        A <= "00010001";
        B <= "00001001";
        C <= "01110101";
        wait for clk_period;
        A <= "11010000";
        B <= "00011100";
        C <= "00000010";
        wait for clk_period;
        A <= "11011110";
        B <= "00110101";
        C <= "11000001";
        wait for clk_period;
        A <= "11101010";
        B <= "01110111";
        C <= "11110010";
        wait for clk_period;
        A <= "11100110";
        B <= "11001010";
        C <= "01111000";
        wait for clk_period;
        A <= "10010000";
        B <= "11100101";
        C <= "11111000";
        wait for clk_period;
        A <= "00100010";
        B <= "00011000";
        C <= "10101010";
        wait for clk_period;
        A <= "01100101";
        B <= "00001111";
        C <= "00101110";
        wait for clk_period;
        A <= "11010100";
        B <= "10010100";
        C <= "00111101";
        wait for clk_period;
        A <= "10011001";
        B <= "00010101";
        C <= "00000011";
        wait for clk_period;
        A <= "00011001";
        B <= "11100111";
        C <= "11101100";
        wait for clk_period;
        A <= "01001101";
        B <= "10010100";
        C <= "01001111";
        wait for clk_period;
        A <= "11111001";
        B <= "01011010";
        C <= "11101010";
        wait for clk_period;
        A <= "10010100";
        B <= "10100010";
        C <= "10001110";
        wait for clk_period;
        A <= "00001100";
        B <= "11001001";
        C <= "01011111";
        wait for clk_period;
        A <= "00000001";
        B <= "01001101";
        C <= "01110110";
        wait for clk_period;
        A <= "01000110";
        B <= "11000001";
        C <= "01101001";
        wait for clk_period;
        A <= "00111011";
        B <= "00001111";
        C <= "10001111";
        wait for clk_period;
        A <= "00001111";
        B <= "01010110";
        C <= "00100110";
        wait for clk_period;
        wait;       
    end process;

end Behavioral;
